* NGSPICE file created from interconnect_inner.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

.subckt interconnect_inner c0_dbg_pc[0] c0_dbg_pc[10] c0_dbg_pc[11] c0_dbg_pc[12]
+ c0_dbg_pc[13] c0_dbg_pc[14] c0_dbg_pc[15] c0_dbg_pc[1] c0_dbg_pc[2] c0_dbg_pc[3]
+ c0_dbg_pc[4] c0_dbg_pc[5] c0_dbg_pc[6] c0_dbg_pc[7] c0_dbg_pc[8] c0_dbg_pc[9] c0_dbg_r0[0]
+ c0_dbg_r0[10] c0_dbg_r0[11] c0_dbg_r0[12] c0_dbg_r0[13] c0_dbg_r0[14] c0_dbg_r0[15]
+ c0_dbg_r0[1] c0_dbg_r0[2] c0_dbg_r0[3] c0_dbg_r0[4] c0_dbg_r0[5] c0_dbg_r0[6] c0_dbg_r0[7]
+ c0_dbg_r0[8] c0_dbg_r0[9] c0_disable c0_i_core_int_sreg[0] c0_i_core_int_sreg[11]
+ c0_i_core_int_sreg[12] c0_i_core_int_sreg[13] c0_i_core_int_sreg[14] c0_i_core_int_sreg[15]
+ c0_i_core_int_sreg[1] c0_i_core_int_sreg[4] c0_i_core_int_sreg[5] c0_i_irq c0_i_mc_core_int
+ c0_i_mem_ack c0_i_mem_data[0] c0_i_mem_data[10] c0_i_mem_data[11] c0_i_mem_data[12]
+ c0_i_mem_data[13] c0_i_mem_data[14] c0_i_mem_data[15] c0_i_mem_data[1] c0_i_mem_data[2]
+ c0_i_mem_data[3] c0_i_mem_data[4] c0_i_mem_data[5] c0_i_mem_data[6] c0_i_mem_data[7]
+ c0_i_mem_data[8] c0_i_mem_data[9] c0_i_mem_exception c0_i_req_data[0] c0_i_req_data[10]
+ c0_i_req_data[11] c0_i_req_data[12] c0_i_req_data[13] c0_i_req_data[14] c0_i_req_data[15]
+ c0_i_req_data[16] c0_i_req_data[17] c0_i_req_data[18] c0_i_req_data[19] c0_i_req_data[1]
+ c0_i_req_data[20] c0_i_req_data[21] c0_i_req_data[22] c0_i_req_data[23] c0_i_req_data[24]
+ c0_i_req_data[25] c0_i_req_data[26] c0_i_req_data[27] c0_i_req_data[28] c0_i_req_data[29]
+ c0_i_req_data[2] c0_i_req_data[30] c0_i_req_data[31] c0_i_req_data[3] c0_i_req_data[4]
+ c0_i_req_data[5] c0_i_req_data[6] c0_i_req_data[7] c0_i_req_data[8] c0_i_req_data[9]
+ c0_i_req_data_valid c0_o_c_data_page c0_o_c_instr_long c0_o_c_instr_page c0_o_icache_flush
+ c0_o_instr_long_addr[0] c0_o_instr_long_addr[1] c0_o_instr_long_addr[2] c0_o_instr_long_addr[3]
+ c0_o_instr_long_addr[4] c0_o_instr_long_addr[5] c0_o_instr_long_addr[6] c0_o_instr_long_addr[7]
+ c0_o_mem_addr[0] c0_o_mem_addr[10] c0_o_mem_addr[11] c0_o_mem_addr[12] c0_o_mem_addr[13]
+ c0_o_mem_addr[14] c0_o_mem_addr[15] c0_o_mem_addr[1] c0_o_mem_addr[2] c0_o_mem_addr[3]
+ c0_o_mem_addr[4] c0_o_mem_addr[5] c0_o_mem_addr[6] c0_o_mem_addr[7] c0_o_mem_addr[8]
+ c0_o_mem_addr[9] c0_o_mem_data[0] c0_o_mem_data[10] c0_o_mem_data[11] c0_o_mem_data[12]
+ c0_o_mem_data[13] c0_o_mem_data[14] c0_o_mem_data[15] c0_o_mem_data[1] c0_o_mem_data[2]
+ c0_o_mem_data[3] c0_o_mem_data[4] c0_o_mem_data[5] c0_o_mem_data[6] c0_o_mem_data[7]
+ c0_o_mem_data[8] c0_o_mem_data[9] c0_o_mem_high_addr[0] c0_o_mem_high_addr[1] c0_o_mem_high_addr[2]
+ c0_o_mem_high_addr[3] c0_o_mem_high_addr[4] c0_o_mem_high_addr[5] c0_o_mem_high_addr[6]
+ c0_o_mem_high_addr[7] c0_o_mem_long_mode c0_o_mem_req c0_o_mem_sel[0] c0_o_mem_sel[1]
+ c0_o_mem_we c0_o_req_active c0_o_req_addr[0] c0_o_req_addr[10] c0_o_req_addr[11]
+ c0_o_req_addr[12] c0_o_req_addr[13] c0_o_req_addr[14] c0_o_req_addr[15] c0_o_req_addr[1]
+ c0_o_req_addr[2] c0_o_req_addr[3] c0_o_req_addr[4] c0_o_req_addr[5] c0_o_req_addr[6]
+ c0_o_req_addr[7] c0_o_req_addr[8] c0_o_req_addr[9] c0_o_req_ppl_submit c0_rst c0_sr_bus_addr[0]
+ c0_sr_bus_addr[10] c0_sr_bus_addr[11] c0_sr_bus_addr[12] c0_sr_bus_addr[13] c0_sr_bus_addr[14]
+ c0_sr_bus_addr[15] c0_sr_bus_addr[1] c0_sr_bus_addr[2] c0_sr_bus_addr[3] c0_sr_bus_addr[4]
+ c0_sr_bus_addr[5] c0_sr_bus_addr[6] c0_sr_bus_addr[7] c0_sr_bus_addr[8] c0_sr_bus_addr[9]
+ c0_sr_bus_data_o[0] c0_sr_bus_data_o[10] c0_sr_bus_data_o[11] c0_sr_bus_data_o[12]
+ c0_sr_bus_data_o[13] c0_sr_bus_data_o[14] c0_sr_bus_data_o[15] c0_sr_bus_data_o[1]
+ c0_sr_bus_data_o[2] c0_sr_bus_data_o[3] c0_sr_bus_data_o[4] c0_sr_bus_data_o[5]
+ c0_sr_bus_data_o[6] c0_sr_bus_data_o[7] c0_sr_bus_data_o[8] c0_sr_bus_data_o[9]
+ c0_sr_bus_we c1_dbg_pc[0] c1_dbg_pc[10] c1_dbg_pc[11] c1_dbg_pc[12] c1_dbg_pc[13]
+ c1_dbg_pc[14] c1_dbg_pc[15] c1_dbg_pc[1] c1_dbg_pc[2] c1_dbg_pc[3] c1_dbg_pc[4]
+ c1_dbg_pc[5] c1_dbg_pc[6] c1_dbg_pc[7] c1_dbg_pc[8] c1_dbg_pc[9] c1_dbg_r0[0] c1_dbg_r0[10]
+ c1_dbg_r0[11] c1_dbg_r0[12] c1_dbg_r0[13] c1_dbg_r0[14] c1_dbg_r0[15] c1_dbg_r0[1]
+ c1_dbg_r0[2] c1_dbg_r0[3] c1_dbg_r0[4] c1_dbg_r0[5] c1_dbg_r0[6] c1_dbg_r0[7] c1_dbg_r0[8]
+ c1_dbg_r0[9] c1_disable c1_i_core_int_sreg[0] c1_i_core_int_sreg[1] c1_i_core_int_sreg[6]
+ c1_i_core_int_sreg[7] c1_i_core_int_sreg[8] c1_i_core_int_sreg[9] c1_i_irq c1_i_mc_core_int
+ c1_i_mem_ack c1_i_mem_data[0] c1_i_mem_data[10] c1_i_mem_data[11] c1_i_mem_data[12]
+ c1_i_mem_data[13] c1_i_mem_data[14] c1_i_mem_data[15] c1_i_mem_data[1] c1_i_mem_data[2]
+ c1_i_mem_data[3] c1_i_mem_data[4] c1_i_mem_data[5] c1_i_mem_data[6] c1_i_mem_data[7]
+ c1_i_mem_data[8] c1_i_mem_data[9] c1_i_mem_exception c1_i_req_data[0] c1_i_req_data[10]
+ c1_i_req_data[11] c1_i_req_data[12] c1_i_req_data[13] c1_i_req_data[14] c1_i_req_data[15]
+ c1_i_req_data[16] c1_i_req_data[17] c1_i_req_data[18] c1_i_req_data[19] c1_i_req_data[1]
+ c1_i_req_data[20] c1_i_req_data[21] c1_i_req_data[22] c1_i_req_data[23] c1_i_req_data[24]
+ c1_i_req_data[25] c1_i_req_data[26] c1_i_req_data[27] c1_i_req_data[28] c1_i_req_data[29]
+ c1_i_req_data[2] c1_i_req_data[30] c1_i_req_data[31] c1_i_req_data[3] c1_i_req_data[4]
+ c1_i_req_data[5] c1_i_req_data[6] c1_i_req_data[7] c1_i_req_data[8] c1_i_req_data[9]
+ c1_i_req_data_valid c1_o_c_data_page c1_o_c_instr_long c1_o_c_instr_page c1_o_icache_flush
+ c1_o_instr_long_addr[0] c1_o_instr_long_addr[1] c1_o_instr_long_addr[2] c1_o_instr_long_addr[3]
+ c1_o_instr_long_addr[4] c1_o_instr_long_addr[5] c1_o_instr_long_addr[6] c1_o_instr_long_addr[7]
+ c1_o_mem_addr[0] c1_o_mem_addr[10] c1_o_mem_addr[11] c1_o_mem_addr[12] c1_o_mem_addr[13]
+ c1_o_mem_addr[14] c1_o_mem_addr[15] c1_o_mem_addr[1] c1_o_mem_addr[2] c1_o_mem_addr[3]
+ c1_o_mem_addr[4] c1_o_mem_addr[5] c1_o_mem_addr[6] c1_o_mem_addr[7] c1_o_mem_addr[8]
+ c1_o_mem_addr[9] c1_o_mem_data[0] c1_o_mem_data[10] c1_o_mem_data[11] c1_o_mem_data[12]
+ c1_o_mem_data[13] c1_o_mem_data[14] c1_o_mem_data[15] c1_o_mem_data[1] c1_o_mem_data[2]
+ c1_o_mem_data[3] c1_o_mem_data[4] c1_o_mem_data[5] c1_o_mem_data[6] c1_o_mem_data[7]
+ c1_o_mem_data[8] c1_o_mem_data[9] c1_o_mem_high_addr[0] c1_o_mem_high_addr[1] c1_o_mem_high_addr[2]
+ c1_o_mem_high_addr[3] c1_o_mem_high_addr[4] c1_o_mem_high_addr[5] c1_o_mem_high_addr[6]
+ c1_o_mem_high_addr[7] c1_o_mem_long_mode c1_o_mem_req c1_o_mem_sel[0] c1_o_mem_sel[1]
+ c1_o_mem_we c1_o_req_active c1_o_req_addr[0] c1_o_req_addr[10] c1_o_req_addr[11]
+ c1_o_req_addr[12] c1_o_req_addr[13] c1_o_req_addr[14] c1_o_req_addr[15] c1_o_req_addr[1]
+ c1_o_req_addr[2] c1_o_req_addr[3] c1_o_req_addr[4] c1_o_req_addr[5] c1_o_req_addr[6]
+ c1_o_req_addr[7] c1_o_req_addr[8] c1_o_req_addr[9] c1_o_req_ppl_submit c1_rst c1_sr_bus_addr[0]
+ c1_sr_bus_addr[10] c1_sr_bus_addr[11] c1_sr_bus_addr[12] c1_sr_bus_addr[13] c1_sr_bus_addr[14]
+ c1_sr_bus_addr[15] c1_sr_bus_addr[1] c1_sr_bus_addr[2] c1_sr_bus_addr[3] c1_sr_bus_addr[4]
+ c1_sr_bus_addr[5] c1_sr_bus_addr[6] c1_sr_bus_addr[7] c1_sr_bus_addr[8] c1_sr_bus_addr[9]
+ c1_sr_bus_data_o[0] c1_sr_bus_data_o[10] c1_sr_bus_data_o[11] c1_sr_bus_data_o[12]
+ c1_sr_bus_data_o[13] c1_sr_bus_data_o[14] c1_sr_bus_data_o[15] c1_sr_bus_data_o[1]
+ c1_sr_bus_data_o[2] c1_sr_bus_data_o[3] c1_sr_bus_data_o[4] c1_sr_bus_data_o[5]
+ c1_sr_bus_data_o[6] c1_sr_bus_data_o[7] c1_sr_bus_data_o[8] c1_sr_bus_data_o[9]
+ c1_sr_bus_we core_clock core_reset dcache_mem_ack dcache_mem_addr[0] dcache_mem_addr[10]
+ dcache_mem_addr[11] dcache_mem_addr[12] dcache_mem_addr[13] dcache_mem_addr[14]
+ dcache_mem_addr[15] dcache_mem_addr[16] dcache_mem_addr[17] dcache_mem_addr[18]
+ dcache_mem_addr[19] dcache_mem_addr[1] dcache_mem_addr[20] dcache_mem_addr[21] dcache_mem_addr[22]
+ dcache_mem_addr[23] dcache_mem_addr[2] dcache_mem_addr[3] dcache_mem_addr[4] dcache_mem_addr[5]
+ dcache_mem_addr[6] dcache_mem_addr[7] dcache_mem_addr[8] dcache_mem_addr[9] dcache_mem_cache_enable
+ dcache_mem_exception dcache_mem_i_data[0] dcache_mem_i_data[10] dcache_mem_i_data[11]
+ dcache_mem_i_data[12] dcache_mem_i_data[13] dcache_mem_i_data[14] dcache_mem_i_data[15]
+ dcache_mem_i_data[1] dcache_mem_i_data[2] dcache_mem_i_data[3] dcache_mem_i_data[4]
+ dcache_mem_i_data[5] dcache_mem_i_data[6] dcache_mem_i_data[7] dcache_mem_i_data[8]
+ dcache_mem_i_data[9] dcache_mem_o_data[0] dcache_mem_o_data[10] dcache_mem_o_data[11]
+ dcache_mem_o_data[12] dcache_mem_o_data[13] dcache_mem_o_data[14] dcache_mem_o_data[15]
+ dcache_mem_o_data[1] dcache_mem_o_data[2] dcache_mem_o_data[3] dcache_mem_o_data[4]
+ dcache_mem_o_data[5] dcache_mem_o_data[6] dcache_mem_o_data[7] dcache_mem_o_data[8]
+ dcache_mem_o_data[9] dcache_mem_req dcache_mem_sel[0] dcache_mem_sel[1] dcache_mem_we
+ dcache_rst dcache_wb_4_burst dcache_wb_ack dcache_wb_adr[0] dcache_wb_adr[10] dcache_wb_adr[11]
+ dcache_wb_adr[12] dcache_wb_adr[13] dcache_wb_adr[14] dcache_wb_adr[15] dcache_wb_adr[16]
+ dcache_wb_adr[17] dcache_wb_adr[18] dcache_wb_adr[19] dcache_wb_adr[1] dcache_wb_adr[20]
+ dcache_wb_adr[21] dcache_wb_adr[22] dcache_wb_adr[23] dcache_wb_adr[2] dcache_wb_adr[3]
+ dcache_wb_adr[4] dcache_wb_adr[5] dcache_wb_adr[6] dcache_wb_adr[7] dcache_wb_adr[8]
+ dcache_wb_adr[9] dcache_wb_cyc dcache_wb_err dcache_wb_i_dat[0] dcache_wb_i_dat[10]
+ dcache_wb_i_dat[11] dcache_wb_i_dat[12] dcache_wb_i_dat[13] dcache_wb_i_dat[14]
+ dcache_wb_i_dat[15] dcache_wb_i_dat[1] dcache_wb_i_dat[2] dcache_wb_i_dat[3] dcache_wb_i_dat[4]
+ dcache_wb_i_dat[5] dcache_wb_i_dat[6] dcache_wb_i_dat[7] dcache_wb_i_dat[8] dcache_wb_i_dat[9]
+ dcache_wb_o_dat[0] dcache_wb_o_dat[10] dcache_wb_o_dat[11] dcache_wb_o_dat[12] dcache_wb_o_dat[13]
+ dcache_wb_o_dat[14] dcache_wb_o_dat[15] dcache_wb_o_dat[1] dcache_wb_o_dat[2] dcache_wb_o_dat[3]
+ dcache_wb_o_dat[4] dcache_wb_o_dat[5] dcache_wb_o_dat[6] dcache_wb_o_dat[7] dcache_wb_o_dat[8]
+ dcache_wb_o_dat[9] dcache_wb_sel[0] dcache_wb_sel[1] dcache_wb_stb dcache_wb_we
+ ic0_mem_ack ic0_mem_addr[0] ic0_mem_addr[10] ic0_mem_addr[11] ic0_mem_addr[12] ic0_mem_addr[13]
+ ic0_mem_addr[14] ic0_mem_addr[15] ic0_mem_addr[1] ic0_mem_addr[2] ic0_mem_addr[3]
+ ic0_mem_addr[4] ic0_mem_addr[5] ic0_mem_addr[6] ic0_mem_addr[7] ic0_mem_addr[8]
+ ic0_mem_addr[9] ic0_mem_cache_flush ic0_mem_data[0] ic0_mem_data[10] ic0_mem_data[11]
+ ic0_mem_data[12] ic0_mem_data[13] ic0_mem_data[14] ic0_mem_data[15] ic0_mem_data[16]
+ ic0_mem_data[17] ic0_mem_data[18] ic0_mem_data[19] ic0_mem_data[1] ic0_mem_data[20]
+ ic0_mem_data[21] ic0_mem_data[22] ic0_mem_data[23] ic0_mem_data[24] ic0_mem_data[25]
+ ic0_mem_data[26] ic0_mem_data[27] ic0_mem_data[28] ic0_mem_data[29] ic0_mem_data[2]
+ ic0_mem_data[30] ic0_mem_data[31] ic0_mem_data[3] ic0_mem_data[4] ic0_mem_data[5]
+ ic0_mem_data[6] ic0_mem_data[7] ic0_mem_data[8] ic0_mem_data[9] ic0_mem_ppl_submit
+ ic0_mem_req ic0_rst ic0_wb_ack ic0_wb_adr[0] ic0_wb_adr[10] ic0_wb_adr[11] ic0_wb_adr[12]
+ ic0_wb_adr[13] ic0_wb_adr[14] ic0_wb_adr[15] ic0_wb_adr[1] ic0_wb_adr[2] ic0_wb_adr[3]
+ ic0_wb_adr[4] ic0_wb_adr[5] ic0_wb_adr[6] ic0_wb_adr[7] ic0_wb_adr[8] ic0_wb_adr[9]
+ ic0_wb_cyc ic0_wb_err ic0_wb_i_dat[0] ic0_wb_i_dat[10] ic0_wb_i_dat[11] ic0_wb_i_dat[12]
+ ic0_wb_i_dat[13] ic0_wb_i_dat[14] ic0_wb_i_dat[15] ic0_wb_i_dat[1] ic0_wb_i_dat[2]
+ ic0_wb_i_dat[3] ic0_wb_i_dat[4] ic0_wb_i_dat[5] ic0_wb_i_dat[6] ic0_wb_i_dat[7]
+ ic0_wb_i_dat[8] ic0_wb_i_dat[9] ic0_wb_sel[0] ic0_wb_sel[1] ic0_wb_stb ic0_wb_we
+ ic1_mem_ack ic1_mem_addr[0] ic1_mem_addr[10] ic1_mem_addr[11] ic1_mem_addr[12] ic1_mem_addr[13]
+ ic1_mem_addr[14] ic1_mem_addr[15] ic1_mem_addr[1] ic1_mem_addr[2] ic1_mem_addr[3]
+ ic1_mem_addr[4] ic1_mem_addr[5] ic1_mem_addr[6] ic1_mem_addr[7] ic1_mem_addr[8]
+ ic1_mem_addr[9] ic1_mem_cache_flush ic1_mem_data[0] ic1_mem_data[10] ic1_mem_data[11]
+ ic1_mem_data[12] ic1_mem_data[13] ic1_mem_data[14] ic1_mem_data[15] ic1_mem_data[16]
+ ic1_mem_data[17] ic1_mem_data[18] ic1_mem_data[19] ic1_mem_data[1] ic1_mem_data[20]
+ ic1_mem_data[21] ic1_mem_data[22] ic1_mem_data[23] ic1_mem_data[24] ic1_mem_data[25]
+ ic1_mem_data[26] ic1_mem_data[27] ic1_mem_data[28] ic1_mem_data[29] ic1_mem_data[2]
+ ic1_mem_data[30] ic1_mem_data[31] ic1_mem_data[3] ic1_mem_data[4] ic1_mem_data[5]
+ ic1_mem_data[6] ic1_mem_data[7] ic1_mem_data[8] ic1_mem_data[9] ic1_mem_ppl_submit
+ ic1_mem_req ic1_rst ic1_wb_ack ic1_wb_adr[0] ic1_wb_adr[10] ic1_wb_adr[11] ic1_wb_adr[12]
+ ic1_wb_adr[13] ic1_wb_adr[14] ic1_wb_adr[15] ic1_wb_adr[1] ic1_wb_adr[2] ic1_wb_adr[3]
+ ic1_wb_adr[4] ic1_wb_adr[5] ic1_wb_adr[6] ic1_wb_adr[7] ic1_wb_adr[8] ic1_wb_adr[9]
+ ic1_wb_cyc ic1_wb_err ic1_wb_i_dat[0] ic1_wb_i_dat[10] ic1_wb_i_dat[11] ic1_wb_i_dat[12]
+ ic1_wb_i_dat[13] ic1_wb_i_dat[14] ic1_wb_i_dat[15] ic1_wb_i_dat[1] ic1_wb_i_dat[2]
+ ic1_wb_i_dat[3] ic1_wb_i_dat[4] ic1_wb_i_dat[5] ic1_wb_i_dat[6] ic1_wb_i_dat[7]
+ ic1_wb_i_dat[8] ic1_wb_i_dat[9] ic1_wb_sel[0] ic1_wb_sel[1] ic1_wb_stb ic1_wb_we
+ inner_disable inner_embed_mode inner_ext_irq inner_wb_4_burst inner_wb_8_burst inner_wb_ack
+ inner_wb_adr[0] inner_wb_adr[10] inner_wb_adr[11] inner_wb_adr[12] inner_wb_adr[13]
+ inner_wb_adr[14] inner_wb_adr[15] inner_wb_adr[16] inner_wb_adr[17] inner_wb_adr[18]
+ inner_wb_adr[19] inner_wb_adr[1] inner_wb_adr[20] inner_wb_adr[21] inner_wb_adr[22]
+ inner_wb_adr[23] inner_wb_adr[2] inner_wb_adr[3] inner_wb_adr[4] inner_wb_adr[5]
+ inner_wb_adr[6] inner_wb_adr[7] inner_wb_adr[8] inner_wb_adr[9] inner_wb_cyc inner_wb_err
+ inner_wb_i_dat[0] inner_wb_i_dat[10] inner_wb_i_dat[11] inner_wb_i_dat[12] inner_wb_i_dat[13]
+ inner_wb_i_dat[14] inner_wb_i_dat[15] inner_wb_i_dat[1] inner_wb_i_dat[2] inner_wb_i_dat[3]
+ inner_wb_i_dat[4] inner_wb_i_dat[5] inner_wb_i_dat[6] inner_wb_i_dat[7] inner_wb_i_dat[8]
+ inner_wb_i_dat[9] inner_wb_o_dat[0] inner_wb_o_dat[10] inner_wb_o_dat[11] inner_wb_o_dat[12]
+ inner_wb_o_dat[13] inner_wb_o_dat[14] inner_wb_o_dat[15] inner_wb_o_dat[1] inner_wb_o_dat[2]
+ inner_wb_o_dat[3] inner_wb_o_dat[4] inner_wb_o_dat[5] inner_wb_o_dat[6] inner_wb_o_dat[7]
+ inner_wb_o_dat[8] inner_wb_o_dat[9] inner_wb_sel[0] inner_wb_sel[1] inner_wb_stb
+ inner_wb_we vccd1 vssd1 c1_i_core_int_sreg[11] c0_i_core_int_sreg[3] c0_i_core_int_sreg[2]
+ c1_i_core_int_sreg[10] c0_i_core_int_sreg[10] c0_i_core_int_sreg[9] c0_i_core_int_sreg[8]
+ c1_i_core_int_sreg[5] c1_i_core_int_sreg[4] c0_i_core_int_sreg[7] c1_i_core_int_sreg[15]
+ c1_i_core_int_sreg[3] c1_i_core_int_sreg[14] c0_i_core_int_sreg[6] c1_i_core_int_sreg[13]
+ c1_i_core_int_sreg[2] c1_i_core_int_sreg[12]
XANTENNA__3140__A1 net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_83_core_clock clknet_3_5_0_core_clock clknet_leaf_83_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3155_ net122 _0905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__3114__I _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3086_ _0845_ net529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6286__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6914_ _0487_ clknet_leaf_57_core_clock dmmu1.page_table\[4\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4640__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input108_I c1_o_c_instr_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6845_ _0418_ clknet_leaf_33_core_clock dmmu0.page_table\[1\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6776_ _0349_ clknet_leaf_100_core_clock dmmu0.long_off_reg\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3988_ net113 immu_1.high_addr_off\[3\] _1650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_9_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5727_ _2758_ _0378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_21_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6145__A1 _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ dmmu0.long_off_reg\[3\] _1803_ _2716_ _2720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input73_I c0_o_req_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4609_ _2059_ _2090_ _2092_ immu_1.page_table\[13\]\[2\] _2095_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5589_ _1976_ _2396_ _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_48_1680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold340 dmmu1.page_table\[5\]\[3\] net1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold351 immu_1.page_table\[5\]\[3\] net1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_2321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4459__A1 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5120__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3131__A1 _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6629__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_2250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5959__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6081__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__CLK clknet_leaf_99_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3895__S _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3198__A1 _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4395__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_2508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3737__A3 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_2519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7166__I net165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6070__I _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6136__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_92_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4870__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4960_ _1817_ _2299_ _2302_ dmmu0.page_table\[7\]\[8\] _2311_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4622__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3911_ _1555_ _1557_ _1301_ _1575_ _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_50_1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ _2264_ _0036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_28_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6630_ _0203_ clknet_leaf_27_core_clock dmmu0.page_table\[12\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6181__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3842_ _1433_ _1507_ _1508_ _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5178__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6561_ _0134_ clknet_leaf_4_core_clock immu_0.page_table\[5\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7076__I net360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3773_ _1410_ _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_55_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5512_ _2637_ _0284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6127__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6492_ _0065_ clknet_leaf_25_core_clock dmmu0.page_table\[14\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5443_ _2596_ _0256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput412 net412 c0_i_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput423 net423 c0_i_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput434 net434 c0_i_req_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5350__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5374_ _2453_ _2553_ _2555_ dmmu0.page_table\[11\]\[2\] _2558_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput445 net445 c0_i_req_data[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput456 net456 c0_i_req_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7113_ net404 net581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3361__A1 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput467 net467 c1_i_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput478 net478 c1_i_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4325_ _1861_ _1911_ _1914_ net949 _1921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput489 net489 c1_i_req_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5638__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7044_ net280 net431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4256_ _1879_ _0595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3207_ _0883_ _0954_ _0940_ _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4187_ _1822_ _0583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input225_I dcache_mem_o_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3138_ _0887_ _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_39_1657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6921__CLK clknet_leaf_64_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_2082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3069_ _0835_ net469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4613__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5810__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6828_ _0401_ clknet_leaf_65_core_clock dmmu1.page_table\[10\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4377__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6759_ _0332_ clknet_leaf_31_core_clock dmmu0.page_table\[5\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6301__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5877__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold170 dmmu0.page_table\[12\]\[8\] net904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_output444_I net444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold181 dmmu1.page_table\[6\]\[6\] net915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold192 dmmu0.page_table\[14\]\[3\] net926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6451__CLK clknet_leaf_23_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4301__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3910__C _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_25_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6109__A1 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3591__A1 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5868__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5332__A2 _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4110_ _1301_ net325 _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_9_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5090_ _2387_ _0112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6944__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4041_ immu_0.page_table\[8\]\[9\] immu_0.page_table\[9\]\[9\] immu_0.page_table\[10\]\[9\]
+ immu_0.page_table\[11\]\[9\] _1463_ _1371_ _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_75_1802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3646__A2 net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4843__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5992_ _2914_ _0487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4943_ _2301_ _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4932__B _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4874_ _1817_ _2242_ _2244_ net837 _2253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6324__CLK clknet_leaf_69_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6613_ _0186_ clknet_leaf_9_core_clock immu_0.page_table\[1\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3825_ immu_0.page_table\[12\]\[3\] immu_0.page_table\[13\]\[3\] _1396_ _1492_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3267__C _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6544_ _0117_ clknet_leaf_18_core_clock immu_0.page_table\[7\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3756_ immu_0.page_table\[4\]\[1\] immu_0.page_table\[5\]\[1\] immu_0.page_table\[12\]\[1\]
+ immu_0.page_table\[13\]\[1\] _1424_ _1377_ _1425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_15_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5571__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6475_ _0048_ clknet_leaf_99_core_clock dmmu0.page_table\[8\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6474__CLK clknet_leaf_10_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3687_ _1348_ net364 _1359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input175_I c1_o_req_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5426_ _2455_ _2582_ _2584_ net824 _2588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_3_984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3334__A1 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4531__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5357_ _2547_ _0219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input342_I ic1_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4308_ _1839_ _1891_ _1909_ _1910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XPHY_EDGE_ROW_58_Left_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5288_ _2507_ _0190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input36_I c0_o_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5087__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4239_ net208 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3637__A2 net260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3193__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_67_Left_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5011__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6817__CLK clknet_leaf_42_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3573__A1 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output659_I net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3325__A1 net150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6967__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Left_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_1734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3420__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4825__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_2020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_2097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6347__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4589__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5250__A1 _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3100__I1 net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3800__A2 _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3239__S1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6497__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3610_ inner_wb_arbiter.o_sel_sig _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5553__A2 _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _2083_ _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_1872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3541_ _1270_ net556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4761__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6260_ _0642_ clknet_leaf_88_core_clock immu_1.page_table\[4\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_2081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5305__A2 _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3472_ _0897_ _1210_ _1211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3316__A1 _1054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5211_ _1811_ _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4513__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6191_ _0573_ clknet_leaf_0_core_clock immu_0.page_table\[11\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5856__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5142_ _2418_ _0133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5069__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _2277_ _2367_ _2369_ net955 _2377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4816__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3619__A2 net266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4024_ net115 immu_1.high_addr_off\[5\] _1684_ _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__3122__I _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ net199 _2889_ _2891_ net744 _2904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ _1837_ _2137_ _2286_ _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_59_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4857_ _2243_ _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_47_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input292_I ic0_mem_data[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_29_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3808_ _1446_ _1475_ _1476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4788_ _1817_ _2191_ _2193_ immu_0.page_table\[12\]\[8\] _2202_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6527_ _0100_ clknet_leaf_7_core_clock immu_0.page_table\[8\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3739_ net366 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_47_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6458_ _0031_ clknet_leaf_23_core_clock dmmu0.page_table\[9\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_2012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3307__A1 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5409_ _2577_ _0241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6389_ _0771_ clknet_leaf_78_core_clock immu_1.page_table\[10\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_2108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3166__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output407_I net407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5232__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3794__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4991__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5535__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7174__I net163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5299__A1 net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_31_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5223__A1 _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3085__I0 net125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5760_ _2777_ _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4711_ _1780_ _2154_ _2155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4982__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5691_ _2738_ _0362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4642_ _2063_ _2108_ _2110_ immu_1.page_table\[12\]\[4\] _2115_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4734__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4573_ _1870_ _2052_ _2054_ immu_1.page_table\[15\]\[10\] _2073_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_2018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6312_ _0694_ clknet_leaf_81_core_clock immu_1.page_table\[3\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3524_ _1261_ net533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6243_ _0625_ clknet_leaf_86_core_clock immu_1.page_table\[2\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3455_ _1193_ _1194_ _0906_ _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3117__I _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6174_ _3018_ _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3386_ net153 dmmu1.long_off_reg\[3\] _1127_ _1128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6512__CLK clknet_leaf_2_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5125_ _2407_ _0127_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3560__I1 net56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input138_I c1_o_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3280__C _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5056_ _2366_ _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4265__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4007_ _1666_ _1667_ _1668_ _1669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__6662__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input305_I ic0_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4017__A2 _1678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5958_ _2895_ _0472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3320__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4909_ _2276_ _0042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5889_ _1873_ _1874_ _2031_ _2855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_75_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5517__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6192__CLK clknet_leaf_1_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3387__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput301 ic0_mem_data[31] net301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput312 ic0_wb_adr[12] net312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output524_I net524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput323 ic0_wb_adr[8] net323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold30 dmmu1.page_table\[9\]\[0\] net764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput334 ic1_mem_data[12] net334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput345 ic1_mem_data[22] net345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold41 immu_1.page_table\[5\]\[6\] net775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput356 ic1_mem_data[3] net356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold52 immu_0.page_table\[4\]\[4\] net786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput367 ic1_wb_adr[13] net367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold63 dmmu0.page_table\[5\]\[0\] net797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput378 ic1_wb_adr[9] net378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold74 dmmu0.page_table\[2\]\[0\] net808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput389 inner_wb_i_dat[0] net389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold85 dmmu0.page_table\[3\]\[7\] net819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_19_1600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold96 dmmu0.page_table\[15\]\[11\] net830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_3_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_97_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_34_core_clock clknet_3_3_0_core_clock clknet_leaf_34_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3697__I _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7169__I net168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3862__S1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3519__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4716__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5417__I _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_5 net390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3365__C _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6535__CLK clknet_leaf_1_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3240_ _0985_ _0986_ _0907_ _0987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5141__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4495__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5692__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3542__I1 net43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3171_ _0889_ _0895_ _0914_ _0920_ _0921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_59_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6685__CLK clknet_leaf_102_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_73_core_clock clknet_3_5_0_core_clock clknet_leaf_73_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_52_1768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5444__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6930_ _0503_ clknet_leaf_55_core_clock dmmu1.page_table\[3\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5995__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _0434_ clknet_leaf_47_core_clock dmmu1.page_table\[8\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7079__I net332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5812_ _2792_ _2802_ _2804_ dmmu1.page_table\[9\]\[6\] _2811_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6792_ _0365_ clknet_leaf_68_core_clock dmmu1.page_table\[13\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3302__S0 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3758__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5743_ _2768_ _0384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3853__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5674_ _2057_ _2726_ _2728_ dmmu1.page_table\[13\]\[1\] _2730_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4625_ _2103_ _2090_ _2092_ immu_1.page_table\[13\]\[9\] _2104_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3275__C _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4556_ _2062_ _0712_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5380__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3507_ _0878_ _1239_ _1244_ _0862_ _1245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_40_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4487_ _1849_ _2014_ _2016_ net901 _2019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input255_I dcache_wb_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6226_ _0608_ clknet_leaf_87_core_clock immu_1.page_table\[0\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3369__S0 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3438_ _0878_ _1175_ _1177_ _1178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4030__S1 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3533__I1 net39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6157_ _1860_ _3000_ _3002_ net940 _3009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3369_ dmmu0.page_table\[8\]\[8\] dmmu0.page_table\[9\]\[8\] dmmu0.page_table\[10\]\[8\]
+ dmmu0.page_table\[11\]\[8\] _0865_ _0868_ _1111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_77_1513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5108_ _1790_ _2396_ _2397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6088_ _2968_ _0529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5039_ _2269_ _2352_ _2354_ immu_0.page_table\[9\]\[3\] _2358_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3997__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6408__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5738__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_2064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4946__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_2583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6163__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_75_2447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_2458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3221__I0 _0967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_75_2469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output641_I net641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5674__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput120 c1_o_mem_addr[11] net120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput131 c1_o_mem_addr[7] net131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput142 c1_o_mem_data[2] net142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput153 c1_o_mem_high_addr[3] net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput164 c1_o_req_addr[0] net164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput175 c1_o_req_addr[5] net175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput186 c1_sr_bus_addr[14] net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4229__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5426__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput197 c1_sr_bus_data_o[0] net197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3421__S _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_2044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5977__A2 _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3988__A1 net113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4401__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4410_ _1969_ _0659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4165__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5390_ _2531_ _2552_ _2554_ dmmu0.page_table\[11\]\[10\] _2566_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput605 net605 ic0_wb_i_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__5901__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput616 net616 ic0_wb_i_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_58_1944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput627 net627 ic1_mem_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4341_ _1846_ _1927_ _1929_ net930 _1931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput638 net638 ic1_mem_req vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_23_996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6179__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput649 net649 ic1_wb_i_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_61_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7060_ net297 net448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_10_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5114__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4272_ _1887_ _0603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6011_ _1770_ _2923_ _2925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3223_ _0955_ _0961_ _0966_ _0970_ net522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__3140__A2 net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3154_ _0897_ _0903_ _0904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3085_ net125 net20 _0842_ _0845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6913_ _0486_ clknet_leaf_52_core_clock dmmu1.page_table\[4\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4640__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6844_ _0417_ clknet_leaf_67_core_clock dmmu1.page_table\[9\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6700__CLK clknet_leaf_35_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3987_ net113 immu_1.high_addr_off\[3\] _1649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6775_ _0348_ clknet_leaf_101_core_clock dmmu0.long_off_reg\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5726_ _2049_ _2742_ _2744_ net1041 _2758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_21_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5657_ _2719_ _0347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6145__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input372_I ic1_wb_adr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6850__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4608_ _2094_ _0732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5588_ _2679_ _0318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input66_I c0_o_req_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3903__A1 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold330 immu_1.page_table\[13\]\[6\] net1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold341 dmmu0.page_table\[15\]\[3\] net1075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4539_ _2049_ _2032_ _2034_ dmmu1.page_table\[14\]\[12\] _2050_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_70_2300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold352 dmmu0.page_table\[1\]\[4\] net1086 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_2322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4459__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6209_ _0591_ clknet_leaf_79_core_clock immu_1.page_table\[9\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7189_ net393 net646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_2240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6230__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5959__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6081__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3514__S0 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6380__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3198__A2 _0939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4395__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_2509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4147__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5344__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5895__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4698__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7182__I net401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_2065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4870__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6723__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4622__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3910_ _1378_ _1560_ _1574_ _1381_ _1575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_80_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4890_ _2258_ _2261_ _2263_ net749 _2264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_28_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3841_ _1474_ immu_1.page_table\[15\]\[3\] _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_15_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6873__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6560_ _0133_ clknet_leaf_6_core_clock immu_0.page_table\[5\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3772_ net366 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_6_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5511_ _2457_ _2630_ _2632_ dmmu0.page_table\[13\]\[4\] _2637_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6491_ _0064_ clknet_leaf_25_core_clock dmmu0.page_table\[14\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6127__A2 _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5442_ _1994_ _2581_ _2583_ net803 _2596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput413 net413 c0_i_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput424 net424 c0_i_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5373_ _2557_ _0225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput435 net435 c0_i_req_data[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_61_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput446 net446 c0_i_req_data[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput457 net457 c0_i_req_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7112_ net403 net580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4324_ _1920_ _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput468 net468 c1_i_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput479 net479 c1_i_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5638__A1 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7043_ net279 net430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4255_ _1824_ _1876_ _1878_ net1006 _1879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6253__CLK clknet_leaf_83_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3206_ _0951_ _0953_ _0878_ _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3744__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4186_ _1821_ _1791_ _1793_ immu_0.page_table\[11\]\[10\] _1822_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3137_ _0886_ _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_37_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input120_I c1_o_mem_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6063__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input218_I dcache_mem_o_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3068_ net216 _0831_ _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5810__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4613__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6827_ _0400_ clknet_leaf_43_core_clock dmmu1.page_table\[10\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3795__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4377__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6758_ _0331_ clknet_leaf_11_core_clock dmmu0.page_table\[6\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5709_ _2749_ _0369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6689_ _0262_ clknet_leaf_90_core_clock immu_1.high_addr_off\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5877__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold160 immu_0.page_table\[5\]\[7\] net894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold171 dmmu0.page_table\[4\]\[6\] net905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold182 dmmu1.page_table\[2\]\[9\] net916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold193 immu_1.page_table\[6\]\[0\] net927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_output437_I net437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4301__A1 net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6746__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_36_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4065__B1 _1718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5652__I1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6896__CLK clknet_leaf_67_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_25_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7177__I net396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5404__I1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5565__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5317__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3591__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__S0 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4040_ immu_0.page_table\[12\]\[9\] immu_0.page_table\[13\]\[9\] immu_0.page_table\[14\]\[9\]
+ immu_0.page_table\[15\]\[9\] _1463_ _1371_ _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_40_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4843__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6045__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _2788_ _2907_ _2909_ dmmu1.page_table\[4\]\[4\] _2914_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_1560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _2300_ _2298_ _2301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_23_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4873_ _2252_ _0030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4359__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6612_ _0185_ clknet_leaf_16_core_clock immu_0.page_table\[1\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3824_ immu_0.page_table\[8\]\[3\] immu_0.page_table\[9\]\[3\] immu_0.page_table\[10\]\[3\]
+ immu_0.page_table\[11\]\[3\] _1370_ _1372_ _1491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_6_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6543_ _0116_ clknet_leaf_19_core_clock immu_0.page_table\[7\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3755_ _1369_ _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_15_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6619__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6474_ _0047_ clknet_leaf_10_core_clock dmmu0.page_table\[8\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3686_ _1356_ _1357_ _1358_ net683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_3_952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_12_Right_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5425_ _2587_ _0247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4531__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5356_ _2527_ _2536_ _2538_ dmmu0.page_table\[15\]\[8\] _2547_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input168_I c1_o_req_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6769__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4307_ _1827_ net181 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
X_5287_ _1802_ _2502_ _2504_ immu_0.page_table\[0\]\[3\] _2507_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5087__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input335_I ic1_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4238_ _1865_ _0591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4295__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input29_I c0_o_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3193__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4169_ _1809_ _1792_ _1794_ immu_0.page_table\[11\]\[5\] _1810_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_21_Right_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5547__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5011__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6299__CLK clknet_leaf_83_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3573__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4770__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Right_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3474__B _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3956__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4286__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4825__A2 _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6027__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4589__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5786__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3649__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3261__A1 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4761__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3540_ net147 net42 _1267_ _1270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6911__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3471_ dmmu1.page_table\[4\]\[11\] dmmu1.page_table\[5\]\[11\] dmmu1.page_table\[6\]\[11\]
+ dmmu1.page_table\[7\]\[11\] _0888_ _0901_ _1210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_10_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5210_ _2460_ _0159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4513__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6190_ _3025_ _3026_ _3027_ _1895_ _0572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4513__B2 dmmu1.page_table\[14\]\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5710__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5141_ _2265_ _2414_ _2416_ immu_0.page_table\[5\]\[1\] _2418_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5072_ _2376_ _0105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4816__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4023_ _1651_ _1682_ _1683_ _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5974_ _2903_ _0480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4925_ net195 net196 _1833_ _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__3252__A1 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6441__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4856_ _1980_ _2241_ _2243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_34_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3807_ immu_1.page_table\[4\]\[2\] immu_1.page_table\[5\]\[2\] immu_1.page_table\[6\]\[2\]
+ immu_1.page_table\[7\]\[2\] _1474_ _1469_ _1475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_15_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4787_ _2201_ _0804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input285_I ic0_mem_data[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6526_ _0099_ clknet_leaf_8_core_clock immu_0.page_table\[8\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3738_ _1407_ _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_31_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6591__CLK clknet_leaf_10_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_2051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6457_ _0030_ clknet_leaf_22_core_clock dmmu0.page_table\[9\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3669_ _1302_ net375 _1345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3307__A2 _1049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5408_ immu_0.high_addr_off\[4\] _1806_ _2572_ _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3938__S0 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6388_ _0770_ clknet_leaf_72_core_clock immu_1.page_table\[10\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5339_ _2537_ _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_60_1968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3166__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6009__A1 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3491__A1 net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_24_core_clock clknet_3_2_0_core_clock clknet_leaf_24_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_70_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5232__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4144__I _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4991__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6934__CLK clknet_leaf_57_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4743__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5299__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7190__I net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_core_clock clknet_3_7_0_core_clock clknet_leaf_63_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6314__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4259__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5471__A2 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_2097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6464__CLK clknet_leaf_23_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4431__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4710_ net85 net84 _2154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4982__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_1547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5690_ _2103_ _2726_ _2728_ net781 _2738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_56_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4641_ _2114_ _0745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4734__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4572_ _2072_ _0718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5931__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6311_ _0693_ clknet_leaf_86_core_clock immu_1.page_table\[3\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3523_ _1246_ _1260_ _0821_ _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6242_ _0624_ clknet_leaf_81_core_clock immu_1.page_table\[2\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3454_ dmmu1.page_table\[0\]\[10\] dmmu1.page_table\[1\]\[10\] dmmu1.page_table\[2\]\[10\]
+ dmmu1.page_table\[3\]\[10\] _0887_ _0909_ _1194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_0_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6173_ dmmu1.long_off_reg\[1\] _1846_ _3016_ _3018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3385_ _1082_ _1125_ _1126_ _1127_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_23_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5124_ _2275_ _2398_ _2400_ immu_0.page_table\[6\]\[6\] _2407_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5055_ _1790_ _2259_ _2366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6807__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4006_ _1666_ _1667_ net2 _1668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4670__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input200_I c1_sr_bus_data_o[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6957__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5957_ _2784_ _2890_ _2892_ net859 _2895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3320__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4908_ _2275_ _2261_ _2263_ net1038 _2276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5888_ _2854_ _0443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input96_I c0_sr_bus_data_o[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4839_ _1812_ _2224_ _2226_ dmmu0.page_table\[10\]\[6\] _2233_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6509_ _0082_ clknet_leaf_109_core_clock immu_0.page_table\[10\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6337__CLK clknet_leaf_71_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4489__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_2386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3387__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3244__S _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput302 ic0_mem_data[3] net302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput313 ic0_wb_adr[13] net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput324 ic0_wb_adr[9] net324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold20 immu_1.page_table\[10\]\[7\] net754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput335 ic1_mem_data[13] net335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold31 dmmu1.page_table\[10\]\[10\] net765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput346 ic1_mem_data[23] net346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold42 immu_1.page_table\[4\]\[2\] net776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput357 ic1_mem_data[4] net357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold53 dmmu1.page_table\[7\]\[9\] net787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6487__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold64 dmmu0.page_table\[5\]\[5\] net798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput368 ic1_wb_adr[14] net368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5989__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput379 ic1_wb_cyc net379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold75 immu_1.page_table\[13\]\[5\] net809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold86 dmmu0.page_table\[12\]\[1\] net820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold97 immu_0.page_table\[13\]\[4\] net831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_19_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4075__S _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_2070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4964__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7185__I net404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4716__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_6 net390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_2030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3662__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5141__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5692__A2 _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3170_ _0915_ _0917_ _0919_ _0920_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_52_1758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5444__A2 _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _0433_ clknet_leaf_47_core_clock dmmu1.page_table\[8\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5811_ _2810_ _0410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3207__A1 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6791_ _0364_ clknet_leaf_40_core_clock dmmu1.page_table\[13\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3302__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5742_ _2065_ _2760_ _2762_ dmmu1.page_table\[11\]\[5\] _2768_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6157__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5673_ _2729_ _0353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_6_Right_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ net209 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_32_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4183__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5380__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4555_ _2061_ _2053_ _2055_ immu_1.page_table\[15\]\[3\] _2062_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3128__I net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3506_ net18 _1241_ _1243_ _1244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_41_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3930__A2 _1582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4486_ _2018_ _0686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6225_ _0607_ clknet_leaf_80_core_clock immu_1.page_table\[0\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5132__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3437_ _0877_ _1176_ _1177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3369__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input150_I c1_o_mem_high_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input248_I dcache_wb_adr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3291__C _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6156_ _3008_ _0557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3368_ dmmu0.page_table\[12\]\[8\] dmmu0.page_table\[13\]\[8\] dmmu0.page_table\[14\]\[8\]
+ dmmu0.page_table\[15\]\[8\] _0865_ _0868_ _1110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3694__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5107_ _2172_ _2296_ _2396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6087_ _2794_ _2958_ _2960_ net872 _2968_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3299_ _0897_ _1043_ _1044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5038_ _2357_ _0090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input11_I c0_o_instr_long_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_2190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6989_ _0562_ clknet_leaf_72_core_clock immu_1.page_table\[8\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_62_2054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4946__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3749__A2 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4422__I _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_2573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_2448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output467_I net467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_2459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output634_I net634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5674__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput110 c1_o_instr_long_addr[0] net110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3685__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput121 c1_o_mem_addr[12] net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_60_1595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput132 c1_o_mem_addr[8] net132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4882__B1 _2243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput143 c1_o_mem_data[3] net143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput154 c1_o_mem_high_addr[4] net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput165 c1_o_req_addr[10] net165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput176 c1_o_req_addr[6] net176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5426__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput187 c1_sr_bus_addr[15] net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput198 c1_sr_bus_data_o[10] net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3437__A1 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4634__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_110_core_clock clknet_3_0_0_core_clock clknet_leaf_110_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_27_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3296__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_45_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6502__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3657__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_59_Right_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3376__C _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_43_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4165__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5362__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput606 net606 ic0_wb_i_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_58_1934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput617 net617 ic0_wb_i_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3912__A2 _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4340_ _1930_ _0628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput628 net628 ic1_mem_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput639 net639 ic1_rst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5114__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4271_ _1866_ _1876_ _1878_ net879 _1887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5163__I _2429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3222_ _0895_ _0969_ _0897_ _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6010_ _2923_ _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_68_Right_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input3_I c0_o_c_instr_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3220__S0 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3153_ dmmu1.page_table\[4\]\[0\] dmmu1.page_table\[5\]\[0\] dmmu1.page_table\[6\]\[0\]
+ dmmu1.page_table\[7\]\[0\] _0899_ _0902_ _0903_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3140__A3 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3084_ _0844_ net518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4625__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6912_ _0485_ clknet_leaf_52_core_clock dmmu1.page_table\[4\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6843_ _0416_ clknet_leaf_42_core_clock dmmu1.page_table\[9\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_1827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4928__A1 net406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6774_ _0347_ clknet_leaf_102_core_clock dmmu0.long_off_reg\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_77_Right_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3986_ _1628_ _1647_ _1648_ net670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5725_ _2757_ _0377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_21_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__I net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input198_I c1_sr_bus_data_o[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5656_ dmmu0.long_off_reg\[2\] _1800_ _2716_ _2719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4607_ _2057_ _2090_ _2092_ immu_1.page_table\[13\]\[1\] _2094_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5587_ _2049_ _2663_ _2665_ dmmu1.page_table\[15\]\[12\] _2679_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold320 immu_0.page_table\[13\]\[7\] net1054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input365_I ic1_wb_adr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold331 dmmu1.page_table\[12\]\[8\] net1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4538_ net200 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xhold342 immu_0.page_table\[14\]\[7\] net1076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold353 dmmu0.page_table\[13\]\[6\] net1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input59_I c0_o_req_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_2323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5105__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4469_ _1860_ _1999_ _2001_ immu_1.page_table\[1\]\[6\] _2008_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_22_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6208_ _0590_ clknet_leaf_73_core_clock immu_1.page_table\[9\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3667__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7188_ net392 net645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4864__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_2007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6139_ _1895_ _2991_ _2997_ _2998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_5_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_2263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3514__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4092__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6525__CLK clknet_leaf_100_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_2016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5041__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output584_I net584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4395__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5592__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4152__I _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6675__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5344__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5895__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_2077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4607__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4083__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3830__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3840_ _1405_ immu_1.page_table\[14\]\[3\] _1507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5583__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3771_ _1439_ _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5510_ _2636_ _0283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6490_ _0063_ clknet_leaf_11_core_clock dmmu0.page_table\[7\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5441_ _2595_ _0255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput414 net414 c0_i_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput425 net425 c0_i_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5372_ _2451_ _2553_ _2555_ dmmu0.page_table\[11\]\[1\] _2557_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3897__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput436 net436 c0_i_req_data[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7111_ net402 net579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput447 net447 c0_i_req_data[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput458 net458 c0_i_req_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4323_ _1858_ _1911_ _1914_ net794 _1920_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput469 net469 c1_i_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5099__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5638__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7042_ net278 net429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4254_ _1877_ _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3649__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3205_ dmmu0.page_table\[12\]\[2\] dmmu0.page_table\[13\]\[2\] dmmu0.page_table\[14\]\[2\]
+ dmmu0.page_table\[15\]\[2\] _0950_ _0952_ _0953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_4185_ net93 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3744__S1 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5621__I _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6548__CLK clknet_leaf_3_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3136_ net120 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_1697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6063__A2 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3067_ _0834_ net468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5271__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input113_I c1_o_instr_long_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5810__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6698__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_1859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6826_ _0399_ clknet_leaf_44_core_clock dmmu1.page_table\[10\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5023__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4377__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6757_ _0330_ clknet_leaf_11_core_clock dmmu0.page_table\[6\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3969_ net8 immu_0.high_addr_off\[3\] _1632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_45_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5708_ _2061_ _2743_ _2745_ net1033 _2749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6688_ _0261_ clknet_leaf_91_core_clock immu_1.high_addr_off\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5639_ _2709_ _0339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5877__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3888__A1 net5 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3432__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold150 dmmu0.page_table\[0\]\[5\] net884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold161 immu_1.page_table\[2\]\[7\] net895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold172 dmmu0.page_table\[9\]\[6\] net906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold183 dmmu1.page_table\[9\]\[10\] net917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold194 immu_1.page_table\[8\]\[5\] net928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4837__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4301__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3499__S0 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3812__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_25_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5565__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3040__A2 net159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5317__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5868__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3879__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3670__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6045__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ _2913_ _0486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6840__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4941_ _1769_ _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_5_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3829__C _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4872_ _1815_ _2242_ _2244_ net974 _2252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6611_ _0184_ clknet_leaf_16_core_clock immu_0.page_table\[1\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6990__CLK clknet_leaf_102_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3823_ _1382_ _1489_ _1378_ _1490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__4006__B net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6542_ _0115_ clknet_leaf_19_core_clock immu_0.page_table\[7\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3754_ immu_0.page_table\[0\]\[1\] immu_0.page_table\[1\]\[1\] immu_0.page_table\[8\]\[1\]
+ immu_0.page_table\[9\]\[1\] _1396_ _1377_ _1423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_27_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6473_ _0046_ clknet_leaf_98_core_clock dmmu0.page_table\[8\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6220__CLK clknet_leaf_84_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3685_ _1337_ net254 _1358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3564__C net533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ _2453_ _2582_ _2584_ net887 _2587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5355_ _2546_ _0218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_7_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4531__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3136__I net120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4306_ _1908_ _0616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5286_ _2506_ _0189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4237_ _1864_ _1841_ _1843_ net1020 _1865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input230_I dcache_wb_4_burst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4295__A1 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input328_I ic0_wb_stb vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4168_ _1808_ _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_14_core_clock clknet_3_2_0_core_clock clknet_leaf_14_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3119_ dmmu0.page_table\[4\]\[0\] dmmu0.page_table\[5\]\[0\] dmmu0.page_table\[6\]\[0\]
+ dmmu0.page_table\[7\]\[0\] _0865_ _0868_ _0869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4047__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4099_ _1535_ net275 _1757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5244__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6809_ _0382_ clknet_leaf_46_core_clock dmmu1.page_table\[11\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5547__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3405__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6713__CLK clknet_leaf_34_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3956__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_53_core_clock clknet_3_7_0_core_clock clknet_leaf_53_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6863__CLK clknet_leaf_48_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5483__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6027__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5786__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7188__I net392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6243__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_92_core_clock clknet_3_4_0_core_clock clknet_leaf_92_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4761__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3470_ _0915_ _1206_ _1208_ _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6393__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4513__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5710__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5140_ _2417_ _0132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5071_ _2275_ _2367_ _2369_ immu_0.page_table\[8\]\[6\] _2376_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3324__I0 _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4022_ net114 immu_1.high_addr_off\[4\] _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4029__A1 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_2070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5973_ _2851_ _2889_ _2891_ net881 _2903_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4924_ _1788_ _2222_ _2284_ _2285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_47_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5529__A1 _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4855_ _2241_ _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_51_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3806_ _1409_ _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_51_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4786_ _1815_ _2191_ _2193_ net911 _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6736__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6525_ _0098_ clknet_leaf_100_core_clock immu_0.page_table\[9\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3737_ net385 _1406_ net107 _1407_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_71_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input180_I c1_o_req_ppl_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3294__C _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input278_I ic0_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6456_ _0029_ clknet_leaf_14_core_clock dmmu0.page_table\[9\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3668_ _1342_ _1343_ _1344_ net679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5407_ _2576_ _0240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3938__S1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ _0769_ clknet_leaf_74_core_clock immu_1.page_table\[10\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6886__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3599_ net213 _1219_ _1300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5338_ _2300_ _2535_ _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input41_I c0_o_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5269_ _1814_ _2486_ _2488_ immu_0.page_table\[1\]\[7\] _2496_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6009__A2 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5217__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6266__CLK clknet_leaf_83_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output497_I net497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4991__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5457__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4743__A2 _2174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4160__I _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_48_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3554__I0 net139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4259__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6609__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5759__A1 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4431__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6759__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4982__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4640_ _2061_ _2108_ _2110_ immu_1.page_table\[12\]\[3\] _2114_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_100_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4734__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ _1868_ _2053_ _2055_ net793 _2072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5931__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6310_ _0692_ clknet_leaf_83_core_clock immu_1.page_table\[3\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3522_ _0894_ _1250_ _1259_ _1260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6241_ _0623_ clknet_leaf_93_core_clock immu_1.page_table\[2\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3453_ dmmu1.page_table\[4\]\[10\] dmmu1.page_table\[5\]\[10\] dmmu1.page_table\[6\]\[10\]
+ dmmu1.page_table\[7\]\[10\] _0887_ _0909_ _1193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4042__S0 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _3017_ _0564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3384_ net152 dmmu1.long_off_reg\[2\] _1126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3170__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5123_ _2406_ _0126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _2365_ _0098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4005_ net9 immu_0.high_addr_off\[4\] _1667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_20_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_50_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4670__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4245__I net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5956_ _2894_ _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4907_ _1811_ _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_63_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5887_ _2049_ _2835_ _2837_ net770 _2854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input395_I inner_wb_i_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4838_ _2232_ _0015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input89_I c0_sr_bus_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4769_ _2190_ _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_16_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6508_ _0081_ clknet_leaf_109_core_clock immu_0.page_table\[10\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6439_ _0012_ clknet_leaf_21_core_clock dmmu0.page_table\[10\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4489__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3525__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3536__I0 net145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5686__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_2387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_4_core_clock clknet_3_0_0_core_clock clknet_leaf_4_core_clock vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_60_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput303 ic0_mem_data[4] net303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold10 dmmu1.page_table\[5\]\[11\] net744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput314 ic0_wb_adr[14] net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold21 immu_1.page_table\[6\]\[9\] net755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput325 net735 net325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_60_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5438__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput336 ic1_mem_data[14] net336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold32 dmmu0.page_table\[0\]\[0\] net766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput347 ic1_mem_data[24] net347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold43 immu_1.page_table\[6\]\[5\] net777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput358 ic1_mem_data[5] net358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5989__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold54 dmmu0.page_table\[5\]\[12\] net788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold65 dmmu0.page_table\[4\]\[5\] net799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput369 ic1_wb_adr[15] net369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold76 dmmu1.page_table\[9\]\[12\] net810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold87 immu_1.page_table\[8\]\[4\] net821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold98 dmmu0.page_table\[14\]\[7\] net832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_3_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6901__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_100_core_clock clknet_3_1_0_core_clock clknet_leaf_100_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4413__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5610__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4964__A2 _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4177__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4716__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5913__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_4_0_core_clock clknet_0_core_clock clknet_3_4_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_7 net391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3527__I0 net141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_2075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5141__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6431__CLK clknet_leaf_108_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4652__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6581__CLK clknet_leaf_4_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _2790_ _2802_ _2804_ dmmu1.page_table\[9\]\[5\] _2810_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6790_ _0363_ clknet_leaf_39_core_clock dmmu1.page_table\[13\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5741_ _2767_ _0383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_2079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5672_ _2051_ _2726_ _2728_ dmmu1.page_table\[13\]\[0\] _2729_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6157__A1 _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4623_ _2102_ _0739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_13_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4554_ _1851_ _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_52_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5380__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3391__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3505_ _0875_ _1242_ _1243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4485_ _1846_ _2014_ _2016_ immu_1.page_table\[3\]\[1\] _2018_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6224_ _0606_ clknet_leaf_82_core_clock immu_1.page_table\[0\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5132__A2 _2397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3436_ dmmu0.page_table\[8\]\[10\] dmmu0.page_table\[9\]\[10\] dmmu0.page_table\[10\]\[10\]
+ dmmu0.page_table\[11\]\[10\] _0871_ _0866_ _1176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3143__A1 net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6155_ _1857_ _3000_ _3002_ net928 _3008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3367_ _1094_ _1109_ net527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input143_I c1_o_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3694__A2 net233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5106_ _2395_ _0120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6086_ _2967_ _0528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6924__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3298_ dmmu1.page_table\[0\]\[5\] dmmu1.page_table\[1\]\[5\] dmmu1.page_table\[2\]\[5\]
+ dmmu1.page_table\[3\]\[5\] _0888_ _0910_ _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_5037_ _2267_ _2352_ _2354_ net961 _2357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input310_I ic0_wb_adr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_2180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6988_ _0561_ clknet_leaf_77_core_clock immu_1.page_table\[8\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4946__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5939_ _2847_ _2873_ _2875_ net959 _2884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_62_2077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6304__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_75_2449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3382__A1 net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6454__CLK clknet_leaf_34_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6171__I1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4331__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3054__I _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput100 c0_sr_bus_data_o[5] net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput111 c1_o_instr_long_addr[1] net111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput122 c1_o_mem_addr[13] net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4882__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3685__A2 net254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput133 c1_o_mem_addr[9] net133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput144 c1_o_mem_data[4] net144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_21_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput155 c1_o_mem_high_addr[5] net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput166 c1_o_req_addr[11] net166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput177 c1_o_req_addr[7] net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput188 c1_sr_bus_addr[1] net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput199 c1_sr_bus_data_o[11] net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_32_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4937__A2 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3296__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6139__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_2115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5362__A2 _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput607 net607 ic0_wb_i_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_58_1935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput618 net618 ic0_wb_i_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_58_1946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput629 net629 ic1_mem_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_58_1957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4270_ _1886_ _0602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5114__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6947__CLK clknet_leaf_64_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3221_ _0967_ _0968_ _0912_ _0969_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_1171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3676__A2 net322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3220__S1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3152_ _0901_ _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3140__A4 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6075__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3083_ net118 net13 _0842_ _0844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3428__A2 _1168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4625__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6911_ _0484_ clknet_leaf_53_core_clock dmmu1.page_table\[4\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6842_ _0415_ clknet_leaf_67_core_clock dmmu1.page_table\[9\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6327__CLK clknet_leaf_61_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6773_ _0346_ clknet_leaf_103_core_clock dmmu0.long_off_reg\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3985_ _1535_ net241 _1648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5724_ _2047_ _2742_ _2744_ dmmu1.page_table\[12\]\[11\] _2757_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5655_ _2718_ _0346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3139__I _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ _2093_ _0731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5586_ _2678_ _0317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3364__A1 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold310 dmmu1.page_table\[15\]\[8\] net1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold321 dmmu1.page_table\[8\]\[4\] net1055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4561__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4537_ _2048_ _0707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold332 dmmu0.page_table\[6\]\[11\] net1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold343 dmmu1.page_table\[5\]\[7\] net1077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input260_I dcache_wb_o_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_2302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_15_Left_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold354 immu_0.page_table\[2\]\[4\] net1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input358_I ic1_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4468_ _2007_ _0679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4313__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6207_ _0589_ clknet_leaf_73_core_clock immu_1.page_table\[9\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3419_ dmmu1.page_table\[12\]\[9\] dmmu1.page_table\[13\]\[9\] dmmu1.page_table\[14\]\[9\]
+ dmmu1.page_table\[15\]\[9\] _0887_ _0900_ _1160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7187_ net391 net644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4399_ _1855_ _1957_ _1959_ net934 _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3667__A2 net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4864__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6138_ _2994_ _0809_ _0810_ _2997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_5_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6069_ _1828_ _1891_ _2030_ _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_68_2242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3602__I _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_2117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A2 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3758__B _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4919__A2 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5041__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5592__A2 _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5465__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5344__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3355__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4552__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3107__A1 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_1810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6057__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4607__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5804__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4083__A2 net245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5280__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3830__A2 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3770_ _1416_ _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_27_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5583__A2 _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5440_ _2531_ _2581_ _2583_ dmmu0.page_table\[2\]\[10\] _2595_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5371_ _2556_ _0224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput415 net415 c0_i_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput426 net426 c0_i_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7110_ net401 net578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput437 net437 c0_i_req_data[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput448 net448 c0_i_req_data[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4322_ _1919_ _0621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput459 net459 c0_i_req_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5099__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7041_ net308 net459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4253_ _1771_ _1875_ _1877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3649__A2 net316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3204_ _0867_ _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4184_ _1820_ _0582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3135_ _0882_ _0883_ _0884_ _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3066_ net215 _0831_ _0834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_54_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5271__A1 net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input106_I c1_o_c_data_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6825_ _0398_ clknet_leaf_49_core_clock dmmu1.page_table\[10\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5023__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3968_ _1581_ _1629_ _1630_ _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_18_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6756_ _0329_ clknet_leaf_11_core_clock dmmu0.page_table\[6\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3585__A1 net229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4782__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5707_ _2748_ _0368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6687_ _0260_ clknet_leaf_91_core_clock immu_1.high_addr_off\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_1002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_2500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3899_ _1463_ immu_0.page_table\[13\]\[5\] _1564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5638_ _1814_ _2699_ _2701_ net1011 _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input71_I c0_o_req_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3337__A1 net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_2034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5569_ _2061_ _2664_ _2666_ dmmu1.page_table\[15\]\[3\] _2670_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3432__S1 _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold140 dmmu0.page_table\[0\]\[9\] net874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold151 immu_1.page_table\[6\]\[1\] net885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold162 dmmu0.page_table\[15\]\[5\] net896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_leaf_43_core_clock clknet_3_6_0_core_clock clknet_leaf_43_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold173 immu_1.page_table\[12\]\[0\] net907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold184 dmmu1.page_table\[2\]\[7\] net918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold195 immu_1.page_table\[12\]\[6\] net929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3533__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4837__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3499__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6642__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_25_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5565__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6792__CLK clknet_leaf_68_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3120__S0 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_82_core_clock clknet_3_5_0_core_clock clknet_leaf_82_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5317__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_105_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4525__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3187__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_55_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4940_ _2298_ _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_75_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4871_ _2251_ _0029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5005__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6610_ _0183_ clknet_leaf_15_core_clock immu_0.page_table\[1\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3822_ _1486_ _1488_ _1366_ _1489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3567__A1 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6541_ _0114_ clknet_leaf_4_core_clock immu_0.page_table\[7\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3753_ icache_arbiter.o_sel_sig _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_42_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6472_ _0045_ clknet_leaf_12_core_clock dmmu0.page_table\[8\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3684_ _1350_ net324 _1326_ _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3319__A1 _1052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5423_ _2586_ _0246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_1339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5354_ _2463_ _2536_ _2538_ dmmu0.page_table\[15\]\[7\] _2546_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_7_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6515__CLK clknet_leaf_8_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4305_ net198 _1893_ _1896_ immu_1.page_table\[0\]\[10\] _1908_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3861__B _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5285_ _1799_ _2502_ _2504_ immu_0.page_table\[0\]\[2\] _2506_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_23_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3178__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4236_ _1863_ _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4295__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4248__I net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_2038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4167_ net100 _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6665__CLK clknet_leaf_104_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3152__I _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input223_I dcache_mem_o_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Left_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3118_ _0867_ _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4098_ _1350_ net329 _1360_ _1756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5244__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3049_ net222 _0822_ _0825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_4_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_2011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6808_ _0381_ clknet_leaf_45_core_clock dmmu1.page_table\[11\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_1455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5547__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4755__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _0312_ clknet_leaf_43_core_clock dmmu1.page_table\[15\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_36_Left_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3405__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6195__CLK clknet_leaf_109_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5180__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output442_I net442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3730__A1 _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4286__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5483__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Left_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_1494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5786__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3797__A1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3341__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4994__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_54_Left_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4621__I net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6538__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_0_core_clock core_clock clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_2084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5710__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6688__CLK clknet_leaf_91_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Left_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5070_ _2375_ _0104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4021_ net114 immu_1.high_addr_off\[4\] _1682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3324__I1 _1065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4029__A2 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5226__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3700__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5972_ _2902_ _0479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3332__S0 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4923_ _1974_ _1782_ _1784_ _2284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_53_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_72_Left_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4854_ _1977_ _2240_ _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_7_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3805_ _1408_ _1472_ _1434_ _1473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_27_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4785_ _2200_ _0803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3736_ net108 _1406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6524_ _0097_ clknet_leaf_2_core_clock immu_0.page_table\[9\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3667_ _1337_ net250 _1344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6455_ _0028_ clknet_leaf_20_core_clock dmmu0.page_table\[9\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3147__I _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_2004 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input173_I c1_o_req_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5406_ immu_0.high_addr_off\[3\] _1803_ _2572_ _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6386_ _0768_ clknet_leaf_78_core_clock immu_1.page_table\[10\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3598_ _1299_ net417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5337_ _2535_ _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3083__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input340_I ic1_mem_data[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5268_ _2495_ _0182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input34_I c0_o_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4219_ net203 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5199_ _1799_ _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6009__A3 _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5217__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3323__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4976__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4728__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3951__A1 net112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6830__CLK clknet_leaf_42_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3554__I1 net34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4259__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6980__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Left_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_50_1698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6210__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5759__A2 _2137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3314__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4431__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6360__CLK clknet_leaf_61_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3395__C _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4570_ _2071_ _0717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5392__B1 _2554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5931__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_2037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3942__A1 net111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3521_ net123 _1253_ _1258_ _0934_ _1259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_53_996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6240_ _0622_ clknet_leaf_86_core_clock immu_1.page_table\[2\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3452_ _1187_ _1190_ _1192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4042__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6171_ dmmu1.long_off_reg\[0\] _1824_ _3016_ _3017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3383_ net152 dmmu1.long_off_reg\[2\] _1125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5122_ _2273_ _2398_ _2400_ net807 _2406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5447__A1 net325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5053_ _2332_ _2351_ _2353_ net828 _2365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4004_ _1631_ _1632_ _1665_ _1666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_46_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4670__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3430__I _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4958__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6703__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5955_ _2782_ _2890_ _2892_ net1091 _2894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _2274_ _0041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5886_ _2853_ _0442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4837_ _1809_ _2224_ _2226_ dmmu0.page_table\[10\]\[5\] _2232_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input290_I ic0_mem_data[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4186__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input388_I inner_wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4768_ _1790_ _2189_ _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6507_ _0080_ clknet_leaf_8_core_clock immu_0.page_table\[10\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3719_ _1370_ immu_0.page_table\[2\]\[0\] _1389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4699_ _2148_ _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6438_ _0011_ clknet_leaf_24_core_clock dmmu0.page_table\[10\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4489__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5686__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3536__I1 net40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_2388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6369_ _0751_ clknet_leaf_77_core_clock immu_1.page_table\[12\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_73_2399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput304 ic0_mem_data[5] net304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3792__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput315 ic0_wb_adr[15] net315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput326 ic0_wb_sel[0] net326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold11 dmmu0.page_table\[9\]\[10\] net745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5438__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold22 dmmu1.page_table\[6\]\[0\] net756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold33 immu_1.page_table\[10\]\[5\] net767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput337 ic1_mem_data[15] net337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput348 ic1_mem_data[25] net348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6233__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold44 dmmu0.page_table\[8\]\[11\] net778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput359 ic1_mem_data[6] net359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold55 dmmu1.page_table\[9\]\[9\] net789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5989__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold66 dmmu1.page_table\[6\]\[7\] net800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4110__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold77 dmmu0.page_table\[3\]\[2\] net811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold88 dmmu0.page_table\[8\]\[3\] net822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold99 dmmu1.page_table\[8\]\[1\] net833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_19_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output405_I net405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_4_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6383__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5610__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4413__A2 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5461__I1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4177__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5374__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_8 net391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_2010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5126__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4101__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6726__CLK clknet_leaf_35_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ _2063_ _2760_ _2762_ net1030 _2767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6876__CLK clknet_leaf_54_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3463__I0 _1186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6157__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5671_ _2727_ _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4622_ _2101_ _2090_ _2092_ net913 _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4553_ _2060_ _0711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3504_ dmmu0.page_table\[12\]\[12\] dmmu0.page_table\[13\]\[12\] dmmu0.page_table\[14\]\[12\]
+ dmmu0.page_table\[15\]\[12\] _0863_ net16 _1242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4484_ _2017_ _0685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5668__A1 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6223_ _0605_ clknet_leaf_92_core_clock immu_1.page_table\[7\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3435_ _0875_ _1174_ _1175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6256__CLK clknet_leaf_93_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6154_ _3007_ _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3774__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3366_ _0860_ _1103_ _1108_ _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_57_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_1505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5105_ _2332_ _2381_ _2383_ immu_0.page_table\[7\]\[10\] _2395_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6085_ _2792_ _2958_ _2960_ net986 _2967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3297_ _0907_ _1041_ _1042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_77_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6093__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input136_I c1_o_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5036_ _2356_ _0089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__A1 _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3160__I _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input303_I ic0_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_2181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6987_ _0560_ clknet_leaf_79_core_clock immu_1.page_table\[8\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_66_2192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5938_ _2883_ _0464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_62_2067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5869_ _2843_ _0435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5356__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_2010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_79_2564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3906__A1 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3536__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3382__A2 net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4331__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput101 c0_sr_bus_data_o[6] net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput112 c1_o_instr_long_addr[2] net112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output522_I net522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput123 c1_o_mem_addr[14] net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4882__A2 _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput134 c1_o_mem_data[0] net134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3271__S _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput145 c1_o_mem_data[5] net145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput156 c1_o_mem_high_addr[6] net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput167 c1_o_req_addr[12] net167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput178 c1_o_req_addr[8] net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput189 c1_sr_bus_addr[2] net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_32_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6899__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3070__A1 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6279__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput608 net608 ic0_wb_i_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_26_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput619 net619 ic0_wb_i_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_58_1947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3220_ dmmu1.page_table\[12\]\[2\] dmmu1.page_table\[13\]\[2\] dmmu1.page_table\[14\]\[2\]
+ dmmu1.page_table\[15\]\[2\] _0889_ _0931_ _0968_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__3756__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3151_ _0900_ _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_20_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6075__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3082_ _0843_ net562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4625__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5822__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6910_ _0483_ clknet_leaf_52_core_clock dmmu1.page_table\[4\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6841_ _0414_ clknet_leaf_65_core_clock dmmu1.page_table\[9\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4389__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6772_ _0345_ clknet_leaf_101_core_clock dmmu0.long_off_reg\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3984_ _1636_ _1646_ _1360_ _1647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5723_ _2756_ _0376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_50_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5654_ dmmu0.long_off_reg\[1\] _1797_ _2716_ _2718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5889__A1 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4605_ _2051_ _2090_ _2092_ net889 _2093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5585_ _2047_ _2663_ _2665_ dmmu1.page_table\[15\]\[11\] _2678_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold300 dmmu0.page_table\[1\]\[10\] net1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4561__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold311 dmmu0.page_table\[8\]\[5\] net1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4536_ _2047_ _2032_ _2034_ net996 _2048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_62_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold322 dmmu0.page_table\[8\]\[7\] net1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_7_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold333 dmmu1.page_table\[6\]\[12\] net1067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_leaf_33_core_clock clknet_3_3_0_core_clock clknet_leaf_33_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold344 dmmu1.page_table\[4\]\[5\] net1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold355 immu_1.page_table\[9\]\[9\] net1089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4467_ _1857_ _1999_ _2001_ immu_1.page_table\[1\]\[5\] _2007_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3155__I net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input253_I dcache_wb_adr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4313__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6206_ _0588_ clknet_leaf_79_core_clock immu_1.page_table\[9\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4313__B2 immu_1.page_table\[2\]\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3747__S0 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3418_ _0894_ _1158_ _1159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4398_ _1963_ _0653_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7186_ net390 net643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4864__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6137_ _2996_ _0550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3349_ _0915_ _1086_ _1091_ _0894_ _1092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_5_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3091__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ _2956_ _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_2243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_2254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5664__I1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5019_ _2275_ _2337_ _2339_ immu_0.page_table\[10\]\[6\] _2346_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5577__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5041__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_72_core_clock clknet_3_4_0_core_clock clknet_leaf_72_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4552__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3107__A2 net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6057__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5804__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3130__I2 _0873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3291__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4624__I net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5656__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4240__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3684__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6914__CLK clknet_leaf_57_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _2444_ _2553_ _2555_ net795 _2556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3977__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput405 net405 c0_disable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput416 net416 c0_i_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput427 net427 c0_i_mem_exception vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput438 net438 c0_i_req_data[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4321_ _1855_ _1911_ _1914_ immu_1.page_table\[2\]\[4\] _1919_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput449 net449 c0_i_req_data[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5099__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4252_ _1875_ _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7040_ net307 net458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3203_ dmmu0.page_table\[4\]\[2\] dmmu0.page_table\[5\]\[2\] dmmu0.page_table\[6\]\[2\]
+ dmmu0.page_table\[7\]\[2\] _0950_ _0948_ _0951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_38_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4183_ _1819_ _1792_ _1794_ immu_0.page_table\[11\]\[9\] _1820_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3134_ _0821_ _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_59_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3065_ _0833_ net482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_1210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5271__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6444__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6824_ _0397_ clknet_leaf_48_core_clock dmmu1.page_table\[10\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5023__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6755_ _0328_ clknet_leaf_37_core_clock dmmu0.page_table\[6\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3967_ net7 immu_0.high_addr_off\[2\] _1630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4782__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3585__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5706_ _2059_ _2743_ _2745_ dmmu1.page_table\[12\]\[2\] _2748_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6686_ _0259_ clknet_leaf_92_core_clock immu_1.high_addr_off\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3898_ _1391_ _1561_ _1562_ _1563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_33_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6594__CLK clknet_leaf_21_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_2501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5637_ _2708_ _0338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input370_I ic1_wb_adr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5568_ _2669_ _0308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input64_I c0_o_req_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold130 dmmu0.page_table\[10\]\[2\] net864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_24_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold141 dmmu0.page_table\[6\]\[9\] net875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_63_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4519_ _1852_ _2033_ _2035_ dmmu1.page_table\[14\]\[3\] _2039_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold152 dmmu1.page_table\[12\]\[5\] net886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5499_ _1976_ _2206_ _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold163 dmmu1.page_table\[13\]\[11\] net897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold174 immu_0.page_table\[10\]\[3\] net908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold185 immu_0.page_table\[15\]\[8\] net919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold196 immu_1.page_table\[5\]\[1\] net930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4837__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7169_ net168 net624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6039__A1 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3273__A1 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3488__C _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6937__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3120__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4525__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4525__B2 dmmu1.page_table\[14\]\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6317__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4289__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3187__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6467__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3264__A1 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4461__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4870_ _1812_ _2242_ _2244_ net906 _2251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3821_ immu_0.page_table\[4\]\[3\] immu_0.page_table\[5\]\[3\] immu_0.page_table\[6\]\[3\]
+ immu_0.page_table\[7\]\[3\] _1487_ _1455_ _1488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__4213__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3567__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6540_ _0113_ clknet_leaf_19_core_clock immu_0.page_table\[7\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3752_ _1308_ _1420_ _1421_ net663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6471_ _0044_ clknet_leaf_22_core_clock dmmu0.page_table\[8\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3683_ _1348_ net378 _1356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5422_ _2451_ _2582_ _2584_ net829 _2586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3319__A2 _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5353_ _2545_ _0217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_7_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4304_ _1907_ _0615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_1529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5284_ _2505_ _0188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3178__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4235_ net207 _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4166_ _1807_ _0577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3117_ _0866_ _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4097_ _1348_ net383 _1755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4047__A3 _1706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5244__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input216_I dcache_mem_o_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3048_ _0824_ net474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_1051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6807_ _0380_ clknet_leaf_47_core_clock dmmu1.page_table\[11\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3809__S _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _1994_ _2316_ _2318_ dmmu0.page_table\[14\]\[11\] _2334_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4755__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_2078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6738_ _0311_ clknet_leaf_43_core_clock dmmu1.page_table\[15\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ _0242_ clknet_leaf_104_core_clock immu_0.high_addr_off\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4507__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5704__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5180__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3544__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output435_I net435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5483__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3494__A1 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output602_I net602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3246__A1 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4994__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3341__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4020_ net659 _1680_ _1681_ net672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5226__A2 _2469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3237__A1 _0982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5971_ _2849_ _2890_ _2892_ dmmu1.page_table\[5\]\[9\] _2902_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_2094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4922_ _2283_ _0048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3332__S1 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4853_ _1779_ _2205_ _2240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_34_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3804_ _1470_ _1471_ _1446_ _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4784_ _1812_ _2191_ _2193_ immu_0.page_table\[12\]\[6\] _2200_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6523_ _0096_ clknet_leaf_2_core_clock immu_0.page_table\[9\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_1697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3735_ _1404_ _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__4033__B _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_2010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _0027_ clknet_leaf_34_core_clock dmmu0.page_table\[9\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3666_ _0814_ net320 _1326_ _1343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5405_ _2575_ _0239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5162__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_2016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6385_ _0767_ clknet_leaf_72_core_clock immu_1.page_table\[10\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6632__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3597_ net220 _1219_ _1299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input166_I c1_o_req_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5336_ _1977_ _2155_ _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_11_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6111__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5267_ _1811_ _2486_ _2488_ immu_0.page_table\[1\]\[6\] _2495_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input333_I ic1_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4218_ _1850_ _0586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3476__A1 net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5198_ _2452_ _0155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6782__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input27_I c0_o_mem_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4149_ _1777_ _1792_ _1794_ immu_0.page_table\[11\]\[0\] _1795_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5217__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4425__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4976__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3323__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4728__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5925__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3400__A1 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5153__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3467__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4664__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3801__I _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3314__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6505__CLK clknet_leaf_3_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5392__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5664__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6655__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3520_ net123 _1255_ _1257_ _1258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_53_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3451_ _1187_ _1190_ _1191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_1359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6170_ _3015_ _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3382_ net1 net53 _1119_ _1123_ _0841_ _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_42_1635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_67_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5121_ _2405_ _0125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5052_ _2364_ _0097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4003_ _1633_ _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4407__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4958__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5954_ _2893_ _0470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4958__B2 dmmu0.page_table\[7\]\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4905_ _2273_ _2261_ _2263_ net1045 _2274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5885_ _2047_ _2835_ _2837_ dmmu1.page_table\[8\]\[11\] _2853_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4836_ _2231_ _0014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5907__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4767_ _1972_ _2154_ _2189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3158__I _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input283_I ic0_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ _0079_ clknet_leaf_0_core_clock immu_0.page_table\[10\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3718_ immu_0.page_table\[1\]\[0\] _1385_ _1387_ _1388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_44_997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4698_ _2065_ _2139_ _2142_ net767 _2148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5135__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6437_ _0010_ clknet_leaf_22_core_clock dmmu0.page_table\[10\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3649_ _0814_ net316 _1326_ _1330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5686__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6368_ _0750_ clknet_leaf_76_core_clock immu_1.page_table\[12\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_2389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5319_ _2461_ _2516_ _2518_ net856 _2525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6299_ _0681_ clknet_leaf_83_core_clock immu_1.page_table\[1\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3792__S1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput305 ic0_mem_data[6] net305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3822__S _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold12 dmmu0.page_table\[5\]\[2\] net746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput316 ic0_wb_adr[1] net316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xinput327 ic0_wb_sel[1] net327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5438__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold23 dmmu0.page_table\[2\]\[9\] net757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput338 ic1_mem_data[16] net338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput349 ic1_mem_data[26] net349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold34 dmmu1.page_table\[3\]\[3\] net768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3449__A1 net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold45 dmmu1.page_table\[6\]\[10\] net779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold56 dmmu1.page_table\[6\]\[3\] net790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4646__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold67 dmmu0.page_table\[6\]\[6\] net801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4110__A2 net325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold78 immu_1.page_table\[15\]\[1\] net812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_58_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold89 dmmu1.page_table\[3\]\[12\] net823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6528__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5071__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5610__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3621__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6678__CLK clknet_leaf_35_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4177__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5374__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_9 net392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5126__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_1955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_1886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4627__I net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4101__A2 net380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5670_ _2682_ _2725_ _2727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_26_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4621_ net208 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_72_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4552_ _2059_ _2053_ _2055_ immu_1.page_table\[15\]\[2\] _2060_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3471__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3503_ _0876_ _1240_ _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_23_core_clock clknet_3_2_0_core_clock clknet_leaf_23_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4483_ _1824_ _2014_ _2016_ immu_1.page_table\[3\]\[0\] _2017_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6222_ _0604_ clknet_leaf_83_core_clock immu_1.page_table\[7\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5668__A2 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3434_ dmmu0.page_table\[12\]\[10\] dmmu0.page_table\[13\]\[10\] dmmu0.page_table\[14\]\[10\]
+ dmmu0.page_table\[15\]\[10\] _0871_ _0866_ _1174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3679__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4876__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6153_ _1854_ _3000_ _3002_ net821 _3007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3774__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3365_ _0860_ _1107_ _0861_ _0821_ _1108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_5104_ _2394_ _0119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6084_ _2966_ _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3296_ dmmu1.page_table\[4\]\[5\] dmmu1.page_table\[5\]\[5\] dmmu1.page_table\[6\]\[5\]
+ dmmu1.page_table\[7\]\[5\] _0888_ _0901_ _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__6093__A2 _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5035_ _2265_ _2352_ _2354_ net972 _2356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input129_I c1_o_mem_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6820__CLK clknet_leaf_48_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6986_ _0559_ clknet_leaf_78_core_clock immu_1.page_table\[8\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_66_2182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5937_ _2794_ _2873_ _2875_ net800 _2883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3603__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3089__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4800__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_2079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_62_core_clock clknet_3_7_0_core_clock clknet_leaf_62_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5868_ _2788_ _2836_ _2838_ net1055 _2843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input94_I c0_sr_bus_data_o[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4819_ _2220_ _0008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6970__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5356__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3206__I1 _0953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3817__S _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5799_ _2803_ _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_79_2565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6200__CLK clknet_leaf_2_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3214__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4331__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3552__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput102 c0_sr_bus_data_o[7] net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput113 c1_o_instr_long_addr[3] net113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput124 c1_o_mem_addr[15] net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6350__CLK clknet_leaf_61_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput135 c1_o_mem_data[10] net135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4619__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput146 c1_o_mem_data[6] net146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_51_1750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput157 c1_o_mem_high_addr[7] net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output515_I net515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput168 c1_o_req_addr[13] net168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4447__I net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput179 c1_o_req_addr[9] net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4095__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3842__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Right_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_1650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4182__I net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3070__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4910__I _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3453__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput609 net609 ic0_wb_i_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_65_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3526__I _1262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Right_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_58_1948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3205__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4858__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3756__S1 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3150_ net121 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6075__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3081_ net162 net57 _0842_ _0843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6843__CLK clknet_leaf_42_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Right_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6840_ _0413_ clknet_leaf_43_core_clock dmmu1.page_table\[9\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5035__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6993__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6771_ _0344_ clknet_leaf_11_core_clock dmmu0.page_table\[5\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5188__I _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3983_ _1348_ _1645_ _1646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5722_ _2105_ _2742_ _2744_ net975 _2756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_1182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5338__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5653_ _2717_ _0345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6223__CLK clknet_leaf_92_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _2091_ _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5889__A2 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5584_ _2677_ _0316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold301 dmmu1.page_table\[10\]\[12\] net1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4535_ net199 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4561__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold312 dmmu0.page_table\[12\]\[10\] net1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold323 dmmu1.page_table\[6\]\[2\] net1057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold334 dmmu1.page_table\[12\]\[7\] net1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold345 immu_0.page_table\[4\]\[9\] net1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold356 immu_0.page_table\[14\]\[3\] net1090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4466_ _2006_ _0678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6373__CLK clknet_leaf_72_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_2315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4849__B1 _2225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6205_ _0587_ clknet_leaf_93_core_clock immu_1.page_table\[9\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4313__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3417_ net154 dmmu1.long_off_reg\[4\] _1157_ _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__3747__S1 _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7185_ net404 net657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4397_ _1852_ _1957_ _1959_ net751 _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input246_I dcache_wb_adr[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6136_ _1771_ _0809_ _0819_ _2995_ _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_22_1869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3348_ _0912_ _1088_ _1090_ _1091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_5_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6067_ net200 _2940_ _2942_ net804 _2956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4077__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Right_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3279_ _0882_ _1023_ _1024_ _0952_ _1025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_68_2244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5018_ _2345_ _0082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_64_2119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5577__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6969_ _0542_ clknet_leaf_58_core_clock dmmu1.page_table\[0\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Right_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4001__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6716__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4552__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output632_I net632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3107__A3 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5501__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6866__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_2069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_73_Right_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_30_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6057__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4068__A1 net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5265__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5804__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3815__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_1605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3130__I3 _0874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5017__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4240__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6396__CLK clknet_leaf_104_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5740__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3977__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput406 net406 c0_i_core_int_sreg[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_65_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput417 net417 c0_i_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4320_ _1918_ _0620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput428 net428 c0_i_req_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput439 net439 c0_i_req_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4251_ _1839_ _1873_ _1874_ _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_43_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3202_ _0864_ _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4182_ net104 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_input1_I c0_o_c_data_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3133_ _0860_ _0861_ _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_21_1880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3064_ net229 _0831_ _0833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_2043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6823_ _0396_ clknet_leaf_48_core_clock dmmu1.page_table\[10\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5559__A1 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6754_ _0327_ clknet_leaf_32_core_clock dmmu0.page_table\[6\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3966_ net7 immu_0.high_addr_off\[2\] _1629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_46_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6739__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5705_ _2747_ _0367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6685_ _0258_ clknet_leaf_102_core_clock icache_arbiter.o_sel_sig vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4782__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3897_ _1385_ immu_0.page_table\[14\]\[5\] _1562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_76_2502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input196_I c1_sr_bus_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5636_ _1811_ _2699_ _2701_ net1048 _2708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5567_ _2059_ _2664_ _2666_ dmmu1.page_table\[15\]\[2\] _2669_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6889__CLK clknet_leaf_54_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input363_I ic1_wb_adr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold120 immu_1.page_table\[11\]\[6\] net854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_14_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4518_ _2038_ _0698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold131 immu_1.page_table\[15\]\[7\] net865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold142 immu_1.page_table\[9\]\[5\] net876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5498_ _2628_ _0279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold153 dmmu0.page_table\[2\]\[2\] net887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input57_I c0_o_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold164 dmmu1.page_table\[2\]\[10\] net898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold175 dmmu1.page_table\[12\]\[6\] net909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold186 immu_1.page_table\[5\]\[7\] net920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4449_ _1995_ _0672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold197 immu_1.page_table\[15\]\[8\] net931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7168_ net167 net623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6039__A2 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6119_ _2847_ _2975_ _2977_ dmmu1.page_table\[0\]\[8\] _2986_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7099_ net354 net507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5798__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6269__CLK clknet_leaf_84_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output582_I net582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4525__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5722__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4289__A1 _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5238__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A1 _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3820_ _1369_ _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4213__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3751_ _1337_ net234 _1421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6470_ _0043_ clknet_leaf_28_core_clock dmmu0.page_table\[8\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3682_ _1353_ _1354_ _1355_ net682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_54_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5421_ _2585_ _0245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5352_ _2461_ _2536_ _2538_ dmmu0.page_table\[15\]\[6\] _2545_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4303_ net209 _1894_ _1897_ immu_1.page_table\[0\]\[9\] _1907_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5283_ _1796_ _2502_ _2504_ immu_0.page_table\[0\]\[1\] _2505_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3714__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5477__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4234_ _1862_ _0590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6411__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4165_ _1806_ _1792_ _1794_ net802 _1807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3116_ net16 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4096_ _1747_ _1753_ _1754_ net675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3047_ net221 _0822_ _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input111_I c1_o_instr_long_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input209_I c1_sr_bus_data_o[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6561__CLK clknet_leaf_4_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6806_ _0379_ clknet_leaf_46_core_clock dmmu1.page_table\[11\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_74_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4998_ _2333_ _0074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4755__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3949_ _1611_ _1612_ net669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6737_ _0310_ clknet_leaf_43_core_clock dmmu1.page_table\[15\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6668_ _0241_ clknet_leaf_103_core_clock immu_0.high_addr_off\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5619_ _2697_ _0331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5704__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6599_ _0172_ clknet_leaf_15_core_clock immu_0.page_table\[2\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3825__S _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5180__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3560__S _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6904__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5640__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4994__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5943__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4190__I net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4054__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_2075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3534__I _1266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6434__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4682__A1 _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6584__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5970_ _2901_ _0478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4921_ _1996_ _2260_ _2262_ dmmu0.page_table\[8\]\[12\] _2283_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4852_ _2239_ _0022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3803_ immu_1.page_table\[0\]\[2\] immu_1.page_table\[1\]\[2\] immu_1.page_table\[2\]\[2\]
+ immu_1.page_table\[3\]\[2\] _1435_ _1469_ _1471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5196__I _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4783_ _2199_ _0802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6522_ _0095_ clknet_leaf_0_core_clock immu_0.page_table\[9\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3734_ net366 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_27_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4033__C net705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6453_ _0026_ clknet_leaf_28_core_clock dmmu0.page_table\[9\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3665_ _1302_ net374 _1342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5404_ immu_0.high_addr_off\[2\] _1800_ _2572_ _2575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3548__I0 net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_2055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6384_ _0766_ clknet_leaf_72_core_clock immu_1.page_table\[10\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3596_ _1298_ net416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5335_ _2534_ _0210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input159_I c1_o_mem_req vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5266_ _2494_ _0181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6111__A1 _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6927__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4217_ _1849_ _1841_ _1843_ net893 _1850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5197_ _2451_ _2447_ _2449_ immu_0.page_table\[3\]\[1\] _2452_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5870__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input326_I ic0_wb_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4148_ _1793_ _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_39_1234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4079_ _1434_ _1738_ _1739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4425__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4976__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6307__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5925__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4728__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6457__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4664__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_2079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4185__I net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3303__B _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6169__A1 _2029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5392__A2 _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_13_core_clock clknet_3_3_0_core_clock clknet_leaf_13_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_52_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3450_ _1157_ _1188_ _1189_ _1190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_46_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3381_ net48 dmmu0.long_off_reg\[3\] _1122_ _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_20_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _2271_ _2398_ _2400_ immu_0.page_table\[6\]\[4\] _2405_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5051_ _2330_ _2352_ _2354_ net818 _2364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4002_ _1422_ _1663_ _1664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3213__B _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4407__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5604__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5953_ _2776_ _2890_ _2892_ net999 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4958__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4904_ _1808_ _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_52_core_clock clknet_3_7_0_core_clock clknet_leaf_52_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5884_ _2852_ _0441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4835_ _1806_ _2224_ _2226_ dmmu0.page_table\[10\]\[4\] _2231_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5907__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4766_ _2188_ _0796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3394__A1 net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6505_ _0078_ clknet_leaf_3_core_clock immu_0.page_table\[10\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3717_ _1386_ _1385_ _1387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4591__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4697_ _2147_ _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input276_I ic0_mem_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6436_ _0009_ clknet_leaf_100_core_clock immu_0.page_table\[13\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3648_ _1302_ net370 _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6183__I1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4343__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6367_ _0749_ clknet_leaf_61_core_clock immu_1.page_table\[12\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3579_ net226 _1204_ _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_60_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5318_ _2524_ _0203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6298_ _0680_ clknet_leaf_87_core_clock immu_1.page_table\[1\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput306 ic0_mem_data[7] net306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput317 ic0_wb_adr[2] net317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xhold13 dmmu1.page_table\[2\]\[0\] net747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput328 ic0_wb_stb net328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xhold24 immu_0.page_table\[6\]\[10\] net758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5249_ _2483_ _0175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput339 ic1_mem_data[17] net339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold35 immu_1.page_table\[7\]\[3\] net769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_23_1591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4646__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold46 dmmu1.page_table\[3\]\[9\] net780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold57 immu_1.page_table\[5\]\[8\] net791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold68 immu_0.page_table\[11\]\[4\] net802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold79 dmmu1.page_table\[10\]\[8\] net813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_leaf_91_core_clock clknet_3_4_0_core_clock clknet_leaf_91_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5071__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3621__A2 net267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output495_I net495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5374__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output662_I net662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4009__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5126__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_2094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3084__I _0844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6087__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5834__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6622__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4620_ _2100_ _0738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3376__A1 _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4551_ _1848_ _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_26_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3502_ dmmu0.page_table\[8\]\[12\] dmmu0.page_table\[9\]\[12\] dmmu0.page_table\[10\]\[12\]
+ dmmu0.page_table\[11\]\[12\] _0863_ net16 _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_40_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3471__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4482_ _2015_ _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_42_2101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6221_ _0603_ clknet_leaf_84_core_clock immu_1.page_table\[7\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4325__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3433_ _1171_ _1172_ _0877_ _1173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5668__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3679__A2 net377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4876__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6152_ _3006_ _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3364_ net47 dmmu0.long_off_reg\[2\] _1106_ _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5103_ _2330_ _2382_ _2384_ immu_0.page_table\[7\]\[9\] _2394_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6083_ _2790_ _2958_ _2960_ net950 _2966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3295_ _1013_ _1040_ net524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__4628__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5034_ _2355_ _0088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_69_Left_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_13_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5053__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6985_ _0558_ clknet_leaf_73_core_clock immu_1.page_table\[8\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_66_2183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5936_ _2882_ _0463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3603__A2 net382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4800__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5867_ _2842_ _0434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input393_I inner_wb_i_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5356__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4818_ _1819_ _2208_ _2210_ immu_0.page_table\[13\]\[9\] _2220_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5798_ _2682_ _2801_ _2803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_7_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input87_I c0_sr_bus_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4564__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4749_ _1800_ _2175_ _2177_ net1032 _2180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6419_ _0801_ clknet_leaf_106_core_clock immu_0.page_table\[12\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3214__S1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput103 c0_sr_bus_data_o[8] net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_60_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput114 c1_o_instr_long_addr[4] net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput125 c1_o_mem_addr[1] net125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_60_1599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7104__I net389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput136 c1_o_mem_data[11] net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4619__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5816__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput147 c1_o_mem_data[7] net147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_51_1751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput158 c1_o_mem_long_mode net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput169 c1_o_req_addr[14] net169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_32_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4095__A2 net246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output508_I net508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6645__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6795__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_45_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4555__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3453__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_0_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3205__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4858__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3080_ _0841_ _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__5283__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_4_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5035__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3982_ _1378_ _1639_ _1644_ _1382_ _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6770_ _0343_ clknet_leaf_38_core_clock dmmu0.page_table\[5\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3597__A1 net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_3_core_clock clknet_3_0_0_core_clock clknet_leaf_3_core_clock vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_35_1281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5721_ _2755_ _0375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_79_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ dmmu0.long_off_reg\[0\] _1777_ _2716_ _2717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5338__A2 _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3349__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4603_ _1912_ _2089_ _2091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4546__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5889__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5583_ _2105_ _2663_ _2665_ dmmu1.page_table\[15\]\[10\] _2677_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4534_ _2046_ _0706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold302 immu_0.page_table\[8\]\[4\] net1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_4_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6518__CLK clknet_leaf_8_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_2430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold313 immu_0.page_table\[13\]\[6\] net1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold324 dmmu1.page_table\[4\]\[7\] net1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold335 immu_0.page_table\[5\]\[4\] net1069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4465_ _1854_ _1999_ _2001_ immu_1.page_table\[1\]\[4\] _2006_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xhold346 dmmu1.page_table\[8\]\[9\] net1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold357 dmmu1.page_table\[5\]\[1\] net1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_2316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4849__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6204_ _0586_ clknet_leaf_93_core_clock immu_1.page_table\[9\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3416_ _1155_ _1127_ _1156_ _1157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7184_ net403 net656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4396_ _1962_ _0652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3521__A1 net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6135_ _2994_ mem_dcache_arb.select _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4548__I _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3347_ _0906_ _1089_ _1090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6668__CLK clknet_leaf_103_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input141_I c1_o_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input239_I dcache_wb_adr[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6066_ _2955_ _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3278_ _0865_ dmmu0.page_table\[0\]\[4\] _1024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_68_2234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5017_ _2273_ _2337_ _2339_ immu_0.page_table\[10\]\[5\] _2345_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_68_2245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5577__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6968_ _0541_ clknet_leaf_57_core_clock dmmu1.page_table\[0\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5919_ _1873_ _1909_ _2031_ _2872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_48_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6899_ _0472_ clknet_leaf_52_core_clock dmmu1.page_table\[5\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6198__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output458_I net458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3107__A4 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5501__A2 _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_81_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3512__A1 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5265__A1 _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3815__A2 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3371__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5017__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3311__B _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3123__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3579__A1 net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4776__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4240__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3537__I _1268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput407 net407 c0_i_core_int_sreg[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_65_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput418 net418 c0_i_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3751__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput429 net429 c0_i_req_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_61_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6810__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4250_ net188 net181 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3201_ _0930_ _0935_ _0947_ _0949_ net521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__4700__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4181_ _1818_ _0581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3132_ _0864_ _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_39_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6960__CLK clknet_leaf_64_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3063_ _0832_ net481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5199__I _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6822_ _0395_ clknet_leaf_46_core_clock dmmu1.page_table\[10\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5559__A2 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6753_ _0326_ clknet_leaf_31_core_clock dmmu0.page_table\[6\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3965_ net107 _1617_ _1627_ _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5704_ _2057_ _2743_ _2745_ dmmu1.page_table\[12\]\[1\] _2747_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3896_ _1463_ immu_0.page_table\[15\]\[5\] _1561_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6684_ _0257_ clknet_leaf_98_core_clock dmmu0.page_table\[2\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6340__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3990__A1 net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4519__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_2503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5635_ _2707_ _0337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input189_I c1_sr_bus_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5566_ _2668_ _0307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold110 immu_1.page_table\[11\]\[3\] net844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold121 dmmu0.page_table\[2\]\[6\] net855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold132 dmmu0.page_table\[13\]\[3\] net866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4517_ _1849_ _2033_ _2035_ dmmu1.page_table\[14\]\[2\] _2038_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5497_ net95 _2612_ _2614_ dmmu0.page_table\[4\]\[12\] _2628_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6490__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold143 immu_1.page_table\[12\]\[7\] net877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold154 dmmu0.page_table\[3\]\[5\] net888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input356_I ic1_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold165 immu_0.page_table\[10\]\[0\] net899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold176 dmmu1.page_table\[4\]\[3\] net910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4448_ _1994_ _1978_ _1981_ dmmu0.page_table\[0\]\[11\] _1995_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold187 dmmu1.page_table\[7\]\[3\] net921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold198 dmmu0.page_table\[13\]\[7\] net932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5495__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4379_ _1864_ _1942_ _1944_ net1050 _1952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7167_ net166 net622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3182__I _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6039__A3 _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6118_ _2985_ _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7098_ net352 net505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_1689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6049_ _2786_ _2941_ _2943_ dmmu1.page_table\[2\]\[3\] _2947_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3558__S _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3981__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6833__CLK clknet_leaf_48_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3733__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4289__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6983__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3092__I _0848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_1955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5238__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3820__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3344__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6363__CLK clknet_leaf_67_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4749__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4213__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3750_ _1401_ _1403_ _1419_ _1350_ _1420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5961__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3681_ _1337_ net253 _1355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5174__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5420_ _2444_ _2582_ _2584_ net808 _2585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3724__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5351_ _2544_ _0216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4302_ _1906_ _0614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5282_ _2500_ _2502_ _2504_ _1386_ _0187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_23_1910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4233_ _1861_ _1841_ _1843_ net1062 _1862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4164_ _1805_ _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_65_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3115_ _0864_ _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4826__I _2225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4095_ _1535_ net246 _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4988__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3046_ _0823_ net467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6706__CLK clknet_leaf_69_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input104_I c0_sr_bus_data_o[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6805_ _0378_ clknet_leaf_68_core_clock dmmu1.page_table\[12\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_1594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ _2332_ _2316_ _2318_ dmmu0.page_table\[14\]\[10\] _2333_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6856__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6736_ _0309_ clknet_leaf_45_core_clock dmmu1.page_table\[15\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3948_ _1306_ net240 _1612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3963__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6667_ _0240_ clknet_leaf_103_core_clock immu_0.high_addr_off\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3879_ _1440_ _1543_ _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5618_ net95 _2680_ _2683_ net753 _2697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4507__A3 _2029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5704__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6598_ _0171_ clknet_leaf_16_core_clock immu_0.page_table\[2\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5549_ _2527_ _2647_ _2649_ dmmu0.page_table\[3\]\[8\] _2658_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_6_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6236__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7112__I net403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6386__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5640__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5943__A2 _2872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3954__A1 net113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_23_Left_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4054__S1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_2065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6729__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4682__A2 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_32_Left_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4920_ _2282_ _0047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6879__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_42_core_clock clknet_3_6_0_core_clock clknet_leaf_42_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_18_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4851_ _1996_ _2223_ _2225_ dmmu0.page_table\[10\]\[12\] _2239_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4198__A1 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3802_ immu_1.page_table\[8\]\[2\] immu_1.page_table\[9\]\[2\] immu_1.page_table\[10\]\[2\]
+ immu_1.page_table\[11\]\[2\] _1435_ _1469_ _1470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_12_1633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4782_ _1809_ _2191_ _2193_ immu_0.page_table\[12\]\[5\] _2199_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3945__A1 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ _0094_ clknet_leaf_3_core_clock immu_0.page_table\[9\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3733_ _0813_ _1402_ _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_55_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_41_Left_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5147__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6452_ _0025_ clknet_leaf_21_core_clock dmmu0.page_table\[9\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3664_ _1339_ _1340_ _1341_ net678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5698__A1 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3548__I1 net31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _2574_ _0238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6259__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3595_ net219 _1219_ _1298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6383_ _0765_ clknet_leaf_74_core_clock immu_1.page_table\[10\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5334_ _1996_ _2515_ _2517_ net784 _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5265_ _1808_ _2486_ _2488_ immu_0.page_table\[1\]\[5\] _2494_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6111__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4122__A1 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4216_ _1848_ _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5196_ _1796_ _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_23_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_50_Left_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5870__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_81_core_clock clknet_3_5_0_core_clock clknet_leaf_81_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4147_ _1771_ _1791_ _1793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_1213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input221_I dcache_mem_o_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3308__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input319_I ic0_wb_adr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4078_ immu_1.page_table\[12\]\[10\] immu_1.page_table\[13\]\[10\] immu_1.page_table\[14\]\[10\]
+ immu_1.page_table\[15\]\[10\] _1404_ _1540_ _1738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5622__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4425__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3029_ mem_dcache_arb.req1_pending net159 _0810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5925__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6719_ _0292_ clknet_leaf_10_core_clock dmmu0.page_table\[13\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7107__I net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_20_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4361__A1 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output440_I net440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput590 net590 ic0_mem_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4113__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__B _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4664__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_2047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_9_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3927__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6401__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3545__I _1272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3380_ _1106_ _1120_ _1121_ _1122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_46_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6551__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5050_ _2363_ _0096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4001_ _1502_ _1657_ _1662_ _1408_ _1663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_20_1946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5852__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5604__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4407__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5455__I1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5952_ _2891_ _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_18_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4903_ _2272_ _0040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5883_ _2851_ _2835_ _2837_ dmmu1.page_table\[8\]\[10\] _2852_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4834_ _2230_ _0013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_1206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5907__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3918__A1 net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4765_ _1821_ _2174_ _2176_ net815 _2188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ _0077_ clknet_leaf_8_core_clock immu_0.page_table\[10\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3716_ net738 _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4591__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4696_ _2063_ _2139_ _2142_ net900 _2147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_1526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6435_ _0008_ clknet_leaf_107_core_clock immu_0.page_table\[13\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3647_ _1325_ _1327_ _1328_ net660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input171_I c1_o_req_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4343__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input269_I dcache_wb_o_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6366_ _0748_ clknet_leaf_75_core_clock immu_1.page_table\[12\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3578_ _1289_ net422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_1835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5317_ _2459_ _2516_ _2518_ net739 _2524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6297_ _0679_ clknet_leaf_86_core_clock immu_1.page_table\[1\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput307 ic0_mem_data[8] net307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold14 dmmu1.page_table\[3\]\[5\] net748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput318 ic0_wb_adr[3] net318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput329 ic0_wb_we net329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5248_ _2332_ _2469_ _2471_ immu_0.page_table\[2\]\[10\] _2483_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input32_I c0_o_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold25 immu_0.page_table\[10\]\[1\] net759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_86_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold36 dmmu1.page_table\[8\]\[12\] net770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4646__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold47 dmmu1.page_table\[13\]\[9\] net781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold58 dmmu0.page_table\[10\]\[10\] net792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold69 dmmu0.page_table\[2\]\[11\] net803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_39_1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5179_ _2439_ _0149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5071__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6424__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3909__A1 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output488_I net488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_7_Left_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6574__CLK clknet_leaf_18_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4009__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4885__A2 _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6087__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5834__A1 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5598__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_2044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6011__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3984__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6917__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3215__I3 dmmu1.page_table\[11\]\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4573__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3376__A2 _1112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4550_ _2058_ _0710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3501_ _1237_ _1238_ _0875_ _1239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4481_ _1912_ _2013_ _2015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6220_ _0602_ clknet_leaf_84_core_clock immu_1.page_table\[7\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4325__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3759__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3432_ dmmu0.page_table\[0\]\[10\] dmmu0.page_table\[1\]\[10\] dmmu0.page_table\[2\]\[10\]
+ dmmu0.page_table\[3\]\[10\] _0871_ _0867_ _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4876__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3363_ _1077_ _1104_ _1105_ _1106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6151_ _1851_ _3000_ _3002_ net740 _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_2380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _2393_ _0118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3294_ net19 _1015_ _1016_ _1039_ _0884_ _1040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6082_ _2965_ _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5033_ _2258_ _2352_ _2354_ net869 _2355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3931__S0 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6447__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6984_ _0557_ clknet_leaf_74_core_clock immu_1.page_table\[8\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_66_2184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5935_ _2792_ _2873_ _2875_ net915 _2882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3064__A1 net229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4261__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4800__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_2095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ _2786_ _2836_ _2838_ net1000 _2842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6597__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4817_ _2219_ _0007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5797_ _2801_ _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_input386_I inner_ext_irq vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4564__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3367__A2 _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4748_ _2179_ _0787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3998__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_2589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4679_ _2135_ _0762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_1_Right_1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5513__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6418_ _0800_ clknet_leaf_104_core_clock immu_0.page_table\[12\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6349_ _0731_ clknet_leaf_60_core_clock immu_1.page_table\[13\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6069__A1 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4010__S _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput104 c0_sr_bus_data_o[9] net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_21_1529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput115 c1_o_instr_long_addr[5] net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput126 c1_o_mem_addr[2] net126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4619__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5816__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput137 c1_o_mem_data[12] net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_1741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput148 c1_o_mem_data[8] net148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_51_1752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput159 c1_o_mem_req net159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_32_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3055__A1 net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4858__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5658__I1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5283__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3294__A1 net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4491__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3294__B2 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7030__I net386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5035__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3981_ _1378_ _1641_ _1643_ _1644_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4243__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5720_ _2103_ _2743_ _2745_ net796 _2755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3597__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5991__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5651_ _2715_ _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4602_ _2089_ _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4546__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3349__A2 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5582_ _2676_ _0315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _1870_ _2032_ _2034_ dmmu1.page_table\[14\]\[10\] _2046_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_74_2420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold303 immu_1.page_table\[6\]\[2\] net1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold314 dmmu0.page_table\[5\]\[6\] net1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold325 dmmu1.page_table\[2\]\[6\] net1059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4464_ _2005_ _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold336 dmmu1.page_table\[0\]\[10\] net1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold347 dmmu1.page_table\[7\]\[1\] net1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4849__A2 _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold358 dmmu0.page_table\[13\]\[9\] net1092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6203_ _0585_ clknet_leaf_80_core_clock immu_1.page_table\[9\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3415_ net153 dmmu1.long_off_reg\[3\] _1156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7183_ net402 net655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4395_ _1849_ _1957_ _1959_ net1037 _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6134_ mem_dcache_arb.transfer_active _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3521__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3346_ dmmu1.page_table\[8\]\[7\] dmmu1.page_table\[9\]\[7\] dmmu1.page_table\[10\]\[7\]
+ dmmu1.page_table\[11\]\[7\] _0898_ _0909_ _1089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6065_ net199 _2940_ _2942_ dmmu1.page_table\[2\]\[11\] _2955_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3277_ dmmu0.page_table\[1\]\[4\] _1023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_input134_I c1_o_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5016_ _2344_ _0081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_68_2246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3285__A1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input301_I ic0_mem_data[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6967_ _0540_ clknet_leaf_55_core_clock dmmu1.page_table\[0\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_2094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5918_ _2871_ _0456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6898_ _0471_ clknet_leaf_53_core_clock dmmu1.page_table\[5\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5849_ _2831_ _0427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5734__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_1738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7115__I net391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6612__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output520_I net520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5265__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4473__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3371__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5017__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4225__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3123__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4776__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3579__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3200__A1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput408 net408 c0_i_irq vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput419 net419 c0_i_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3751__A2 net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3553__I _1276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3200_ _0948_ _0862_ _0842_ _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4700__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4180_ _1817_ _1792_ _1794_ immu_0.page_table\[11\]\[8\] _1818_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_1603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3131_ _0862_ _0880_ _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3062_ net228 _0831_ _0832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3267__A1 net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3267__B2 _1012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_2110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6821_ _0394_ clknet_leaf_47_core_clock dmmu1.page_table\[10\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5559__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4767__A1 _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6752_ _0325_ clknet_leaf_13_core_clock dmmu0.page_table\[6\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3964_ _0813_ _1626_ _1627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5703_ _2746_ _0366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6683_ _0256_ clknet_leaf_98_core_clock dmmu0.page_table\[2\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3895_ _1558_ _1559_ _1367_ _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4519__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5634_ _1808_ _2699_ _2701_ net798 _2707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4519__B2 dmmu1.page_table\[14\]\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5716__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5192__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5565_ _2057_ _2664_ _2666_ net1022 _2668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6635__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold100 dmmu0.page_table\[2\]\[8\] net834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_14_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold111 immu_1.page_table\[3\]\[9\] net845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4516_ _2037_ _0697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_1315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold122 dmmu0.page_table\[12\]\[6\] net856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold133 immu_1.page_table\[3\]\[4\] net867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5496_ _2627_ _0278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_1949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold144 immu_0.page_table\[4\]\[10\] net878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold155 immu_1.page_table\[13\]\[0\] net889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold166 immu_1.page_table\[10\]\[4\] net900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4447_ net94 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xhold177 immu_0.page_table\[12\]\[7\] net911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input251_I dcache_wb_adr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold188 dmmu1.page_table\[10\]\[2\] net922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_25_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold199 immu_1.page_table\[5\]\[2\] net933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5495__A2 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input349_I ic1_mem_data[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7166_ net165 net621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4378_ _1951_ _0645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6785__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6117_ _1863_ _2975_ _2977_ dmmu1.page_table\[0\]\[7\] _2985_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3329_ dmmu0.page_table\[0\]\[6\] dmmu0.page_table\[1\]\[6\] dmmu0.page_table\[2\]\[6\]
+ dmmu0.page_table\[3\]\[6\] _0872_ _0941_ _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7097_ net351 net504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6048_ _2946_ _0511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3258__A1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3839__S _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5955__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4930__A1 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4694__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4997__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3344__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_32_core_clock clknet_3_3_0_core_clock clknet_leaf_32_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6508__CLK clknet_leaf_109_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4749__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6658__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3680_ _1350_ net323 _1326_ _1354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5174__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5350_ _2459_ _2536_ _2538_ net896 _2544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4921__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4301_ net208 _1894_ _1897_ immu_1.page_table\[0\]\[8\] _1906_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5281_ _2503_ _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5477__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_2093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4232_ _1860_ _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3488__A1 _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_71_core_clock clknet_3_4_0_core_clock clknet_leaf_71_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4163_ net99 _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3114_ _0863_ _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4094_ _1750_ _1751_ _1752_ _1360_ _1753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_21_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4437__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3232__B _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4988__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3045_ net214 _0822_ _0823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6804_ _0377_ clknet_leaf_40_core_clock dmmu1.page_table\[12\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5937__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4996_ net93 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_19_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_2086 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6735_ _0308_ clknet_leaf_45_core_clock dmmu1.page_table\[15\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3947_ net659 _1594_ _1610_ _1611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_19_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3412__A1 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6666_ _0239_ clknet_leaf_104_core_clock immu_0.high_addr_off\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input299_I ic0_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3963__A2 _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3878_ immu_1.page_table\[8\]\[5\] immu_1.page_table\[9\]\[5\] immu_1.page_table\[10\]\[5\]
+ immu_1.page_table\[11\]\[5\] _1404_ _1540_ _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5617_ _2696_ _0330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6597_ _0170_ clknet_leaf_19_core_clock immu_0.page_table\[2\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5548_ _2657_ _0300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input62_I c0_o_req_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5479_ _2455_ _2613_ _2615_ net997 _2619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_6_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4676__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7149_ net404 net619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_1498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_2016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_93_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6105__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6330__CLK clknet_leaf_71_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_2086 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5758__I _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6480__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4850_ _2238_ _0021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_1650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3801_ _1410_ _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_51_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4781_ _2198_ _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6520_ _0093_ clknet_leaf_109_core_clock immu_0.page_table\[9\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3732_ _1370_ _1382_ _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5147__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6451_ _0024_ clknet_leaf_23_core_clock dmmu0.page_table\[9\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3663_ _1337_ net249 _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5402_ immu_0.high_addr_off\[1\] _1797_ _2572_ _2574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5698__A2 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6382_ _0764_ clknet_leaf_78_core_clock immu_1.page_table\[10\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3594_ _1297_ net415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3227__B _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5333_ _2533_ _0209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5264_ _2493_ _0180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4215_ net202 _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4122__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5195_ _2450_ _0154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5870__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4146_ _1791_ _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3881__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3308__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6823__CLK clknet_leaf_48_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4077_ _1440_ _1736_ _1737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input214_I dcache_mem_o_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5622__A2 _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3028_ mem_dcache_arb.req0_pending net54 _0809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3633__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3389__S _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6973__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4979_ _2322_ _0066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6718_ _0291_ clknet_leaf_12_core_clock dmmu0.page_table\[13\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6649_ _0222_ clknet_leaf_12_core_clock dmmu0.page_table\[15\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6203__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4361__A2 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6353__CLK clknet_leaf_61_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput580 net580 dcache_wb_i_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput591 net591 ic0_mem_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_output433_I net433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7123__I net68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1004 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_1075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5301__A1 net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3561__I _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7033__I net288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4000_ _1415_ _1659_ _1661_ _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5852__A2 _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3863__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5065__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5604__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ _1770_ _2889_ _2891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3615__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6996__CLK clknet_leaf_95_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4812__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4902_ _2271_ _2261_ _2263_ net902 _2272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5882_ net198 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_34_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5368__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4833_ _1803_ _2224_ _2226_ net1052 _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6226__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4764_ _2187_ _0795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6503_ _0076_ clknet_leaf_9_core_clock dmmu0.page_table\[14\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3715_ _1384_ _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_70_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4591__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4695_ _2146_ _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6434_ _0007_ clknet_leaf_107_core_clock immu_0.page_table\[13\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3646_ _1306_ net231 _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6376__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4343__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6365_ _0747_ clknet_leaf_75_core_clock immu_1.page_table\[12\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3577_ net225 _1204_ _1289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_45_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input164_I c1_o_req_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5316_ _2523_ _0202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6296_ _0678_ clknet_leaf_81_core_clock immu_1.page_table\[1\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput308 ic0_mem_data[9] net308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5247_ _2482_ _0174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput319 ic0_wb_adr[4] net319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xhold15 dmmu0.page_table\[8\]\[0\] net749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold26 immu_0.page_table\[4\]\[1\] net760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input331_I ic1_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold37 immu_0.page_table\[5\]\[8\] net771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold48 dmmu1.page_table\[10\]\[9\] net782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold59 immu_1.page_table\[15\]\[9\] net793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5178_ _2275_ _2430_ _2432_ immu_0.page_table\[4\]\[6\] _2439_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input25_I c0_o_mem_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _1775_ net658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_3_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3606__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3847__S _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4031__A1 _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6719__CLK clknet_leaf_10_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__I net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5531__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6869__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6087__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4098__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5834__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3845__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5047__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_2012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5598__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6249__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3757__S _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4940__I _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6011__A2 _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4022__A1 net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6399__CLK clknet_leaf_108_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3456__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3500_ dmmu0.page_table\[4\]\[12\] dmmu0.page_table\[5\]\[12\] dmmu0.page_table\[6\]\[12\]
+ dmmu0.page_table\[7\]\[12\] _0863_ _0866_ _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_48_1847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4480_ _2013_ _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3208__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4325__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3431_ dmmu0.page_table\[4\]\[10\] dmmu0.page_table\[5\]\[10\] dmmu0.page_table\[6\]\[10\]
+ dmmu0.page_table\[7\]\[10\] _0871_ _0867_ _1171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3759__S1 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5771__I _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6150_ _3005_ _0554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3362_ net46 dmmu0.long_off_reg\[1\] _1105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_72_2370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _2328_ _2382_ _2384_ immu_0.page_table\[7\]\[8\] _2393_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6081_ _2788_ _2958_ _2960_ net982 _2965_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4089__A1 net116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3293_ _0879_ _1021_ _1026_ _1031_ _1038_ _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_77_1509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5032_ _2353_ _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3836__A1 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3931__S1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5589__A1 _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6983_ _0556_ clknet_leaf_79_core_clock immu_1.page_table\[8\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_1520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_66_2174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_2185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5934_ _2881_ _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_2196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4261__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3064__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5865_ _2841_ _0433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4816_ _1817_ _2208_ _2210_ immu_0.page_table\[13\]\[8\] _2219_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5796_ _1829_ _2031_ _2801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_69_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4747_ _1797_ _2175_ _2177_ net890 _2179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4564__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5761__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3998__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input281_I ic0_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input379_I ic1_wb_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4678_ _2103_ _2123_ _2125_ net1005 _2135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6417_ _0799_ clknet_leaf_106_core_clock immu_0.page_table\[12\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5513__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3629_ _0812_ net271 _1318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6348_ _0730_ clknet_leaf_70_core_clock immu_1.page_table\[14\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6069__A2 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput105 c0_sr_bus_we net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6279_ _0661_ clknet_leaf_33_core_clock dmmu0.page_table\[0\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput116 c1_o_instr_long_addr[6] net116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput127 c1_o_mem_addr[3] net127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_51_1731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5816__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput138 c1_o_mem_data[13] net138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_1742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput149 c1_o_mem_data[9] net149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_51_1753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3827__A1 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3055__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6541__CLK clknet_leaf_4_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_32_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4555__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5752__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6691__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5591__I _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4491__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3980_ _1368_ _1642_ _1643_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4243__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5440__B1 _2583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4794__A2 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5991__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5650_ _1975_ _2570_ _2715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _1828_ _1839_ _2028_ _2089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_5_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4546__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5581_ _2103_ _2664_ _2666_ net936 _2676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4532_ _2045_ _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_2421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold304 dmmu0.page_table\[8\]\[6\] net1038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold315 dmmu0.page_table\[4\]\[7\] net1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_2443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4463_ _1851_ _1999_ _2001_ immu_1.page_table\[1\]\[3\] _2005_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xhold326 immu_1.page_table\[13\]\[10\] net1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold337 immu_1.page_table\[5\]\[5\] net1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold348 dmmu1.page_table\[1\]\[8\] net1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_61_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_2307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6202_ _0584_ clknet_leaf_79_core_clock immu_1.page_table\[9\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3414_ net153 dmmu1.long_off_reg\[3\] _1155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_70_2318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_15_Right_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7182_ net401 net654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4394_ _1961_ _0651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6133_ _1771_ _0810_ _0822_ _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_26_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3345_ _0896_ _1087_ _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6414__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5259__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6064_ _2954_ _0519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3276_ dmmu0.page_table\[2\]\[4\] dmmu0.page_table\[3\]\[4\] _0865_ _1022_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5015_ _2271_ _2337_ _2339_ immu_0.page_table\[10\]\[4\] _2344_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_2236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_2247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3285__A2 _1027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input127_I c1_o_mem_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6564__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Right_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6966_ _0539_ clknet_leaf_57_core_clock dmmu1.page_table\[0\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5917_ _2049_ _2855_ _2857_ dmmu1.page_table\[7\]\[12\] _2871_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6897_ _0470_ clknet_leaf_52_core_clock dmmu1.page_table\[5\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _2529_ _2819_ _2821_ dmmu0.page_table\[1\]\[9\] _2831_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input92_I c0_sr_bus_data_o[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5734__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5779_ _2791_ _0397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_98_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_33_Right_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3145__B _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_10_Left_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output513_I net513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7131__I net61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4473__A1 net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_22_core_clock clknet_3_2_0_core_clock clknet_leaf_22_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_73_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Right_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3028__A2 net54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4225__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5422__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4776__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3100__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_51_Right_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3200__A2 _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput409 net409 c0_i_mc_core_int vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6437__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5489__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4161__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4700__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_61_core_clock clknet_3_7_0_core_clock clknet_leaf_61_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3130_ _0869_ _0870_ _0873_ _0874_ _0877_ _0879_ _0880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6587__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3061_ _0821_ _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_59_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7041__I net308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_60_Right_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_2100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _0393_ clknet_leaf_48_core_clock dmmu1.page_table\[10\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_2111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_2011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6751_ _0324_ clknet_leaf_30_core_clock dmmu0.page_table\[6\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3963_ _1502_ _1620_ _1625_ _1408_ _1626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_58_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5702_ _2051_ _2743_ _2745_ net987 _2746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6682_ _0255_ clknet_leaf_97_core_clock dmmu0.page_table\[2\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3894_ immu_0.page_table\[0\]\[5\] immu_0.page_table\[1\]\[5\] immu_0.page_table\[2\]\[5\]
+ immu_0.page_table\[3\]\[5\] _1487_ _1390_ _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4519__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5716__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ _2706_ _0336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5564_ _2667_ _0306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4515_ _1846_ _2033_ _2035_ dmmu1.page_table\[14\]\[1\] _2037_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold101 dmmu0.page_table\[8\]\[2\] net835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold112 immu_0.page_table\[14\]\[4\] net846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold123 dmmu1.page_table\[10\]\[5\] net857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5495_ net94 _2612_ _2614_ dmmu0.page_table\[4\]\[11\] _2627_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold134 dmmu1.page_table\[1\]\[9\] net868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold145 immu_1.page_table\[7\]\[8\] net879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold156 immu_0.page_table\[14\]\[1\] net890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4446_ _1993_ _0671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6141__A1 _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold167 immu_1.page_table\[3\]\[2\] net901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold178 dmmu1.page_table\[1\]\[2\] net912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_10_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold189 immu_1.page_table\[10\]\[0\] net923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7165_ net179 net635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4377_ _1861_ _1942_ _1944_ net991 _1951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_1625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input244_I dcache_wb_adr[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6116_ _2984_ _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3328_ dmmu0.page_table\[4\]\[6\] dmmu0.page_table\[5\]\[6\] dmmu0.page_table\[6\]\[6\]
+ dmmu0.page_table\[7\]\[6\] _0872_ _0941_ _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7096_ net350 net503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6047_ _2784_ _2941_ _2943_ dmmu1.page_table\[2\]\[2\] _2946_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3259_ dmmu1.page_table\[15\]\[4\] _1005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4455__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3412__C _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5400__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4207__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5955__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _0522_ clknet_leaf_53_core_clock dmmu1.page_table\[1\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_25_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3855__S _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3194__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4391__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7126__I net71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6132__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output630_I net630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4694__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4997__A2 _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4749__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5174__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3185__A1 net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7036__I net303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4921__A2 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4300_ _1905_ _0613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5280_ _1895_ _2501_ _2503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6123__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4231_ net206 _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_23_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4162_ _1804_ _0576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3113_ net15 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4093_ _1748_ _1731_ _1749_ _1752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4437__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5634__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3044_ _0821_ _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4988__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6803_ _0376_ clknet_leaf_68_core_clock dmmu1.page_table\[12\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5937__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__I net366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4995_ _2331_ _0073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6734_ _0307_ clknet_leaf_44_core_clock dmmu1.page_table\[15\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3946_ _1422_ _1605_ _1609_ _1610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_30_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3412__A2 _1147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6665_ _0238_ clknet_leaf_104_core_clock immu_0.high_addr_off\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3877_ _1434_ _1541_ _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input194_I c1_sr_bus_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5616_ net94 _2680_ _2683_ net1066 _2696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6596_ _0169_ clknet_leaf_5_core_clock immu_0.page_table\[2\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4373__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6752__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5547_ _2463_ _2647_ _2649_ net819 _2657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input361_I ic1_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5478_ _2618_ _0269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_1769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input55_I c0_o_mem_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4429_ _1800_ _1979_ _1982_ dmmu0.page_table\[0\]\[2\] _1985_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_1460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3479__A2 _1214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7148_ net403 net618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7079_ net332 net485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_1518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6282__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_1961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3167__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6105__A1 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6625__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5919__A1 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3559__I _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3800_ _1383_ _1460_ _1467_ _1468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_12_1613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4780_ _1806_ _2191_ _2193_ net805 _2198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3731_ _1374_ _1379_ _1382_ _1400_ _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_51_1695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5774__I _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3662_ _0814_ net319 _1326_ _1340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5147__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6450_ _0023_ clknet_leaf_22_core_clock dmmu0.page_table\[9\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5401_ _2573_ _0237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4355__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6381_ _0763_ clknet_leaf_72_core_clock immu_1.page_table\[11\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5698__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3593_ net218 _1219_ _1297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_45_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ _1994_ _2515_ _2517_ dmmu0.page_table\[12\]\[11\] _2533_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_51_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_2069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5263_ _1805_ _2486_ _2488_ immu_0.page_table\[1\]\[4\] _2493_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4658__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4214_ _1847_ _0585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5194_ _2444_ _2447_ _2449_ immu_0.page_table\[3\]\[0\] _2450_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4145_ _1781_ _1790_ _1791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_78_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4076_ immu_1.page_table\[8\]\[10\] immu_1.page_table\[9\]\[10\] immu_1.page_table\[10\]\[10\]
+ immu_1.page_table\[11\]\[10\] _1404_ _1540_ _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_78_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5083__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3633__A2 net258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input207_I c1_sr_bus_data_o[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4978_ _2267_ _2317_ _2319_ net952 _2322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3397__A1 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6717_ _0290_ clknet_leaf_12_core_clock dmmu0.page_table\[13\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_1934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3929_ _1382_ _1587_ _1592_ _1593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA_clkbuf_leaf_37_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6648_ _0221_ clknet_leaf_10_core_clock dmmu0.page_table\[15\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6579_ _0152_ clknet_leaf_3_core_clock immu_0.page_table\[4\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4361__A3 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput570 net570 dcache_wb_i_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput581 net581 dcache_wb_i_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5846__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput592 net592 ic0_mem_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_57_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6648__CLK clknet_leaf_10_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6798__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6023__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4585__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6177__I1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4888__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5950_ _2889_ _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_18_1833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4812__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3615__A2 net264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4901_ _1805_ _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_73_1172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ _2850_ _0440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4832_ _2229_ _0012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5368__A2 _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3379__A1 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4763_ _1819_ _2175_ _2177_ immu_0.page_table\[14\]\[9\] _2187_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _0075_ clknet_leaf_13_core_clock dmmu0.page_table\[14\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3714_ _1369_ _1384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4694_ _2061_ _2139_ _2142_ net962 _2146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6433_ _0006_ clknet_leaf_106_core_clock immu_0.page_table\[13\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3645_ _0814_ net309 _1326_ _1327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3576_ _1288_ net421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6364_ _0746_ clknet_leaf_77_core_clock immu_1.page_table\[12\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5315_ _2457_ _2516_ _2518_ dmmu0.page_table\[12\]\[4\] _2523_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6295_ _0677_ clknet_leaf_88_core_clock immu_1.page_table\[1\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input157_I c1_o_mem_high_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput309 ic0_wb_adr[0] net309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5246_ _2330_ _2470_ _2472_ net1053 _2482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold16 dmmu1.page_table\[10\]\[11\] net750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold27 immu_1.page_table\[7\]\[6\] net761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3303__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold38 dmmu1.page_table\[13\]\[6\] net772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold49 dmmu0.page_table\[12\]\[9\] net783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5177_ _2438_ _0148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input324_I ic0_wb_adr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4128_ _0812_ net230 _1775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_39_1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6940__CLK clknet_leaf_57_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I c0_o_mem_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4059_ immu_0.page_table\[8\]\[10\] immu_0.page_table\[9\]\[10\] immu_0.page_table\[10\]\[10\]
+ immu_0.page_table\[11\]\[10\] _1487_ _1390_ _1719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_36_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3606__A2 net328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3199__I _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4567__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6320__CLK clknet_leaf_69_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4319__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5531__A2 _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7134__I net64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6470__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4098__A2 net329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__A1 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3845__A2 _1511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5047__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5598__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3153__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4558__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3456__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3081__I0 net162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_13_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3781__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3208__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3430_ _1170_ net530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3361_ net46 dmmu0.long_off_reg\[1\] _1104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4730__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7044__I net280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_29_Left_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5100_ _2392_ _0117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_72_2382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6080_ _2964_ _0525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3292_ _0938_ _1034_ _1037_ _0878_ _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__6963__CLK clknet_leaf_54_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5031_ _2140_ _2351_ _2353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3392__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6982_ _0555_ clknet_leaf_73_core_clock immu_1.page_table\[8\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_2175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5933_ _2790_ _2873_ _2875_ dmmu1.page_table\[6\]\[5\] _2881_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_66_2186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_2197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4261__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5864_ _2784_ _2836_ _2838_ net1072 _2841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_2097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6343__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4549__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4815_ _2218_ _0006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5795_ _2800_ _0404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4746_ _2178_ _0786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_2569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6493__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4677_ _2134_ _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input274_I dcache_wb_stb vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6416_ _0798_ clknet_leaf_105_core_clock immu_0.page_table\[12\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5513__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3628_ _1317_ net699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6347_ _0729_ clknet_leaf_76_core_clock immu_1.page_table\[14\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3559_ _1279_ net560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6069__A3 _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6278_ _0660_ clknet_leaf_92_core_clock immu_1.page_table\[6\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput106 c1_o_c_data_page net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput117 c1_o_instr_long_addr[7] net117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput128 c1_o_mem_addr[4] net128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_51_1732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput139 c1_o_mem_data[14] net139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5229_ _2473_ _0165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_51_1743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_12_core_clock clknet_3_3_0_core_clock clknet_leaf_12_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5202__I _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_1672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output493_I net493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7129__I net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_2085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6836__CLK clknet_leaf_48_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3763__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4960__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6986__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3606__B net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_51_core_clock clknet_3_7_0_core_clock clknet_leaf_51_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6216__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4491__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6366__CLK clknet_leaf_75_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4243__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5440__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5991__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_2050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7039__I net306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4600_ _2088_ _0730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5580_ _2675_ _0314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_90_core_clock clknet_3_4_0_core_clock clknet_leaf_90_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _1868_ _2033_ _2035_ dmmu1.page_table\[14\]\[9\] _2045_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_2422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold305 immu_0.page_table\[4\]\[3\] net1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold316 immu_1.page_table\[4\]\[7\] net1050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_68_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4462_ _2004_ _0676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold327 immu_1.page_table\[14\]\[6\] net1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold338 dmmu1.page_table\[8\]\[2\] net1072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold349 dmmu0.page_table\[13\]\[2\] net1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_7_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6201_ _0583_ clknet_leaf_100_core_clock immu_0.page_table\[11\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3506__A1 net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_2308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3413_ _1144_ _1153_ _0840_ _1154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_26_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_2319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4393_ _1846_ _1957_ _1959_ net885 _1961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_1954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7181_ net400 net653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6132_ _1771_ _2992_ _2993_ _0548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_26_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3344_ dmmu1.page_table\[12\]\[7\] dmmu1.page_table\[13\]\[7\] dmmu1.page_table\[14\]\[7\]
+ dmmu1.page_table\[15\]\[7\] _0887_ _0909_ _1087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_0_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5259__A1 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3275_ _0948_ _1017_ _1020_ _0877_ _1021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_42_1299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6063_ _2851_ _2940_ _2942_ net898 _2954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5014_ _2343_ _0080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6709__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_2248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6965_ _0538_ clknet_leaf_51_core_clock dmmu1.page_table\[0\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6859__CLK clknet_leaf_48_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5916_ _2870_ _0455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_2069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6896_ _0469_ clknet_leaf_67_core_clock dmmu1.page_table\[6\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5847_ _2830_ _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input391_I inner_wb_i_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5778_ _2790_ _2778_ _2780_ net857 _2791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5734__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input85_I c0_sr_bus_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4729_ _2166_ _0781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3426__B net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6239__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3356__S0 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6389__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4473__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5670__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output506_I net506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_47_1609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4225__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5422__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A2 _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3984__A1 _1636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4933__B1 _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5489__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4161__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3060_ _0830_ net480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_1903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_2047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_63_2101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5777__I _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6750_ _0323_ clknet_leaf_28_core_clock dmmu0.page_table\[6\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3962_ _1415_ _1622_ _1624_ _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_57_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5701_ _2744_ _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_72_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6681_ _0254_ clknet_leaf_38_core_clock dmmu0.page_table\[2\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3893_ immu_0.page_table\[4\]\[5\] immu_0.page_table\[5\]\[5\] immu_0.page_table\[6\]\[5\]
+ immu_0.page_table\[7\]\[5\] _1487_ _1455_ _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_6_913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5632_ _1805_ _2699_ _2701_ dmmu0.page_table\[5\]\[4\] _2706_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5716__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3727__A1 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5563_ _2051_ _2664_ _2666_ dmmu1.page_table\[15\]\[0\] _2667_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4514_ _2036_ _0696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold102 immu_0.page_table\[2\]\[5\] net836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold113 dmmu1.page_table\[8\]\[5\] net847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5494_ _2626_ _0277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold124 dmmu1.page_table\[3\]\[10\] net858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold135 immu_0.page_table\[9\]\[0\] net869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold146 immu_1.page_table\[4\]\[1\] net880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4445_ _1821_ _1978_ _1981_ dmmu0.page_table\[0\]\[10\] _1993_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold157 immu_0.page_table\[10\]\[7\] net891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6141__A2 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold168 dmmu0.page_table\[8\]\[4\] net902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold179 immu_1.page_table\[13\]\[8\] net913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7164_ net178 net634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4376_ _1950_ _0644_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6531__CLK clknet_leaf_109_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6115_ _1860_ _2975_ _2977_ dmmu1.page_table\[0\]\[6\] _2984_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_1659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3327_ _0934_ _1068_ _1070_ _1051_ _0841_ _1071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7095_ net349 net502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input237_I dcache_wb_adr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5101__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6046_ _2945_ _0510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3258_ _0931_ _1000_ _1003_ _0897_ _1004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_55_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3189_ _0877_ _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6681__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input404_I inner_wb_i_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6948_ _0521_ clknet_leaf_63_core_clock dmmu1.page_table\[2\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5955__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3966__A1 net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6879_ _0452_ clknet_leaf_59_core_clock dmmu1.page_table\[7\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5168__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4915__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4391__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4930__A3 _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output456_I net456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4143__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5340__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_2_core_clock clknet_3_0_0_core_clock clknet_leaf_2_core_clock vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_9_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4694__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5891__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_109_core_clock clknet_3_0_0_core_clock clknet_leaf_109_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7142__I net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3329__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_44_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6404__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3709__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6554__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6123__A2 _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4134__A1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4230_ _1859_ _0589_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4161_ _1803_ _1792_ _1794_ immu_0.page_table\[11\]\[3\] _1804_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7052__I net289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3112_ _0860_ _0861_ _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4092_ _0813_ net107 _1751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5634__A1 _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4437__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3043_ _0819_ _0820_ _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_72_1023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6802_ _0375_ clknet_leaf_66_core_clock dmmu1.page_table\[12\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4994_ _2330_ _2317_ _2319_ dmmu0.page_table\[14\]\[9\] _2331_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5937__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3948__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6733_ _0306_ clknet_leaf_45_core_clock dmmu1.page_table\[15\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3945_ net107 _1608_ _1609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6664_ _0237_ clknet_leaf_104_core_clock immu_0.high_addr_off\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3876_ immu_1.page_table\[12\]\[5\] immu_1.page_table\[13\]\[5\] immu_1.page_table\[14\]\[5\]
+ immu_1.page_table\[15\]\[5\] _1404_ _1540_ _1541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5615_ _2695_ _0329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3755__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6595_ _0168_ clknet_leaf_21_core_clock immu_0.page_table\[2\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4373__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input187_I c1_sr_bus_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5546_ _2656_ _0299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5477_ _2453_ _2613_ _2615_ dmmu0.page_table\[4\]\[2\] _2618_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_1136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input354_I ic1_mem_data[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4428_ _1984_ _0662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_6_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input48_I c0_o_mem_high_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7147_ net402 net617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4359_ _1870_ _1926_ _1928_ net1025 _1940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7078_ net362 net515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6029_ _2847_ _2924_ _2926_ net925 _2935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6427__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4027__S _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3939__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_1804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6577__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5400__I1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_2079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6105__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5313__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5864__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_0_0_core_clock clknet_0_core_clock clknet_3_0_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_79_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5616__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_2011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5467__I1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5919__A2 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6041__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3776__S _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3730_ _1383_ _1393_ _1399_ _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_3_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3661_ _1302_ net373 _1339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7047__I net283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5400_ immu_0.high_addr_off\[0\] _1777_ _2572_ _2573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4355__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3789__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6380_ _0762_ clknet_leaf_77_core_clock immu_1.page_table\[11\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3592_ _1296_ net414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5331_ _2532_ _0208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4107__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5262_ _2492_ _0179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4213_ _1846_ _1841_ _1843_ immu_1.page_table\[9\]\[1\] _1847_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5193_ _2448_ _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4144_ _1789_ _1790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_39_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4075_ _1733_ _1734_ _1439_ _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4291__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input102_I c0_sr_bus_data_o[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4977_ _2321_ _0065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6716_ _0289_ clknet_leaf_13_core_clock dmmu0.page_table\[13\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3397__A2 net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3928_ _1378_ _1589_ _1591_ _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_62_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6647_ _0220_ clknet_leaf_13_core_clock dmmu0.page_table\[15\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3859_ _1368_ _1524_ _1525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_1979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5543__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6578_ _0151_ clknet_leaf_18_core_clock immu_0.page_table\[4\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5529_ _1976_ _2445_ _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__5406__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6099__A1 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput560 net560 dcache_mem_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput571 net571 dcache_wb_i_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5846__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput582 net582 ic0_mem_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput593 net593 ic0_mem_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_79_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5205__I _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6023__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4585__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4337__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4888__A2 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3076__A1 net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6742__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4273__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4812__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4900_ _2270_ _0039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5880_ _2849_ _2836_ _2838_ net1080 _2850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_1184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4831_ _1800_ _2224_ _2226_ net864 _2229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_56_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6892__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _2186_ _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6501_ _0074_ clknet_leaf_10_core_clock dmmu0.page_table\[14\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3713_ _1377_ _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_55_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4693_ _2145_ _0766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6432_ _0005_ clknet_leaf_108_core_clock immu_0.page_table\[13\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3644_ _1304_ _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5525__B1 _2631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6363_ _0745_ clknet_leaf_67_core_clock immu_1.page_table\[12\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3575_ net224 _1204_ _1288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_23_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5314_ _2522_ _0201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6294_ _0676_ clknet_leaf_87_core_clock immu_1.page_table\[1\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5828__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6272__CLK clknet_leaf_84_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5245_ _2481_ _0173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold17 immu_1.page_table\[6\]\[3\] net751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold28 immu_1.page_table\[11\]\[7\] net762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_23_1595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5176_ _2273_ _2430_ _2432_ immu_0.page_table\[4\]\[5\] _2438_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold39 dmmu0.page_table\[9\]\[2\] net773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_39_1002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4127_ net659 _0816_ net565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_58_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input317_I ic0_wb_adr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4058_ _1383_ _1715_ _1717_ _1718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_56_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6005__A1 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_1989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4319__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_41_core_clock clknet_3_6_0_core_clock clknet_leaf_41_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3164__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6765__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7150__I net390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5047__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4255__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3153__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4558__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_80_core_clock clknet_3_5_0_core_clock clknet_leaf_80_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5507__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6295__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4730__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3360_ _1096_ _1098_ _1100_ _1102_ _1103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_42_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_2361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3291_ _0882_ _1035_ _1036_ _0948_ _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_5030_ _2351_ _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3297__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3392__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3049__A1 net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3521__C _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6981_ _0554_ clknet_leaf_73_core_clock immu_1.page_table\[8\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5932_ _2880_ _0461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_66_2176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_1653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_2187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5863_ _2840_ _0432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4814_ _1815_ _2208_ _2210_ net1054 _2218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4549__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5746__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5794_ _2049_ _2777_ _2779_ net1035 _2800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4745_ _1777_ _2175_ _2177_ net946 _2178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6638__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4676_ _2101_ _2123_ _2125_ immu_1.page_table\[11\]\[8\] _2134_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6415_ _0797_ clknet_leaf_106_core_clock immu_0.page_table\[12\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3627_ _1308_ net270 _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input267_I dcache_wb_o_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6346_ _0728_ clknet_leaf_75_core_clock immu_1.page_table\[14\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3558_ net160 net55 _0841_ _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6788__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6277_ _0659_ clknet_leaf_83_core_clock immu_1.page_table\[6\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3489_ net50 dmmu0.long_off_reg\[5\] _1228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput107 c1_o_c_instr_long net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput118 c1_o_mem_addr[0] net118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5228_ _2444_ _2470_ _2472_ immu_0.page_table\[2\]\[0\] _2473_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3288__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput129 c1_o_mem_addr[5] net129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_51_1733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input30_I c0_o_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4485__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5159_ _2332_ _2413_ _2415_ immu_0.page_table\[5\]\[10\] _2427_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_32_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_49_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4237__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4788__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5985__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_2020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3460__A1 net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output486_I net486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3212__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3874__S _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4960__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3673__I _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7145__I net400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3279__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_101_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5440__A2 _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_2040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_51_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ _2044_ _0704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6930__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_2423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold306 immu_0.page_table\[12\]\[0\] net1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4461_ _1848_ _1999_ _2001_ immu_1.page_table\[1\]\[2\] _2004_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6153__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_2434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold317 immu_1.page_table\[7\]\[1\] net1051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold328 immu_1.page_table\[9\]\[6\] net1062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6200_ _0582_ clknet_leaf_2_core_clock immu_0.page_table\[11\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold339 immu_0.page_table\[7\]\[5\] net1073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3412_ _0878_ _1147_ _1152_ _0883_ _1153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_7180_ net399 net652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_70_2309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4392_ _1960_ _0650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6131_ net559 _2991_ mem_dcache_arb.select _2993_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3343_ _1084_ _1085_ _0896_ _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_1868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5259__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6062_ _2953_ _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3274_ _0882_ _1018_ _1019_ _0952_ _1020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4467__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5013_ _2269_ _2337_ _2339_ net908 _2343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_2238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__CLK clknet_leaf_83_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3690__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5967__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3817__I0 net236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6964_ _0537_ clknet_leaf_56_core_clock dmmu1.page_table\[0\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_2086 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5915_ _2047_ _2855_ _2857_ dmmu1.page_table\[7\]\[11\] _2870_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3442__A1 net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6895_ _0468_ clknet_leaf_65_core_clock dmmu1.page_table\[6\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6460__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5846_ _2527_ _2819_ _2821_ dmmu0.page_table\[1\]\[8\] _2830_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5777_ _1857_ _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_20_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input384_I inner_disable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4728_ _1812_ _2157_ _2159_ immu_0.page_table\[15\]\[6\] _2166_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4942__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input78_I c0_sr_bus_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4659_ _2124_ _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_32_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_1920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_2019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6329_ _0711_ clknet_leaf_74_core_clock immu_1.page_table\[15\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5414__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3356__S1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_5_0_core_clock clknet_0_core_clock clknet_3_5_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5670__A2 _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_48_Left_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3681__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6803__CLK clknet_leaf_68_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5422__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5186__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6953__CLK clknet_leaf_57_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Left_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4933__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4933__B2 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5489__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4161__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6333__CLK clknet_leaf_71_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5110__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Left_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_1038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6483__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3961_ _1440_ _1623_ _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5700_ _2682_ _2742_ _2744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_70_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6680_ _0253_ clknet_leaf_37_core_clock dmmu0.page_table\[2\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3892_ net2 _1556_ _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_75_Left_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5631_ _2705_ _0335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5562_ _2665_ _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_14_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4513_ _1824_ _2033_ _2035_ dmmu1.page_table\[14\]\[0\] _2036_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5493_ _2531_ _2612_ _2614_ dmmu0.page_table\[4\]\[10\] _2626_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold103 dmmu0.page_table\[9\]\[8\] net837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold114 immu_1.page_table\[2\]\[2\] net848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold125 dmmu1.page_table\[5\]\[2\] net859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold136 immu_0.page_table\[3\]\[9\] net870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4444_ _1992_ _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold147 dmmu1.page_table\[5\]\[10\] net881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4688__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold158 immu_0.page_table\[3\]\[10\] net892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6141__A3 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold169 dmmu0.page_table\[6\]\[2\] net903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7163_ net177 net633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4375_ _1858_ _1942_ _1944_ immu_1.page_table\[4\]\[5\] _1950_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3360__B1 _1100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6114_ _2983_ _0540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3326_ net151 dmmu1.long_off_reg\[1\] _1069_ _1070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7094_ net348 net501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_2074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6045_ _2782_ _2941_ _2943_ net942 _2945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_2085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5101__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3257_ _0889_ _1001_ _1002_ _0902_ _1003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__6826__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input132_I c1_o_mem_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3663__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3188_ dmmu0.page_table\[8\]\[1\] dmmu0.page_table\[9\]\[1\] dmmu0.page_table\[10\]\[1\]
+ dmmu0.page_table\[11\]\[1\] _0872_ _0868_ _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4860__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6976__CLK clknet_leaf_102_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3415__A1 net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6947_ _0520_ clknet_leaf_64_core_clock dmmu1.page_table\[2\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6878_ _0451_ clknet_leaf_55_core_clock dmmu1.page_table\[7\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5168__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5829_ _2820_ _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6206__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3718__A2 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4915__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6117__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4391__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5208__I _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6356__CLK clknet_leaf_61_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5340__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output449_I net449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3741__I2 immu_1.page_table\[2\]\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3329__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3654__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__B1 _2225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3900__B _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4134__A2 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6849__CLK clknet_leaf_34_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4160_ _1802_ _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_65_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3111_ net1 net53 _0861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_65_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4091_ _1748_ _1731_ _1749_ _1750_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_21_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5095__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5634__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3042_ mem_dcache_arb.select net559 _0820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6999__CLK clknet_leaf_103_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput290 ic0_mem_data[21] net290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3645__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6801_ _0374_ clknet_leaf_42_core_clock dmmu1.page_table\[12\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4993_ net104 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_59_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6229__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_2007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3101__I _0853_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3944_ net112 immu_1.high_addr_off\[2\] _1607_ _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__3948__A2 net240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6732_ _0305_ clknet_leaf_98_core_clock dmmu0.page_table\[3\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6663_ _0236_ clknet_leaf_100_core_clock dmmu0.page_table\[11\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3875_ _1410_ _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_45_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5614_ _2531_ _2680_ _2683_ dmmu0.page_table\[6\]\[10\] _2695_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6379__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6594_ _0167_ clknet_leaf_21_core_clock immu_0.page_table\[2\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_1197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4373__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5545_ _2461_ _2647_ _2649_ net969 _2656_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5476_ _2617_ _0268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4427_ _1797_ _1979_ _1982_ dmmu0.page_table\[0\]\[1\] _1984_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3771__I _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input347_I ic1_mem_data[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7146_ net401 net616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4358_ _1939_ _0637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3309_ _0938_ _1053_ _1054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7077_ net361 net514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4289_ _1848_ _1894_ _1897_ immu_1.page_table\[0\]\[2\] _1900_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_59_2070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6028_ _2934_ _0503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4833__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5561__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5313__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7153__I net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5077__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5616__A2 _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3627__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6041__A2 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3486__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6521__CLK clknet_leaf_3_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3660_ _1335_ _1336_ _1338_ net677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3238__S0 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4355__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3591_ net217 _1219_ _1296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3789__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5330_ _2531_ _2515_ _2517_ net1046 _2532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3805__B _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4107__A2 net273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5261_ _1802_ _2486_ _2488_ immu_0.page_table\[1\]\[3\] _2492_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_45_1479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4212_ _1845_ _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_62_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5192_ _1980_ _2446_ _2448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4143_ _1769_ _1785_ _1788_ _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_23_1788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4074_ immu_1.page_table\[0\]\[10\] immu_1.page_table\[1\]\[10\] immu_1.page_table\[2\]\[10\]
+ immu_1.page_table\[3\]\[10\] _1435_ _1469_ _1734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_74_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4291__A1 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4976_ _2265_ _2317_ _2319_ net994 _2321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_1237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5240__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6715_ _0288_ clknet_leaf_23_core_clock dmmu0.page_table\[13\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3766__I _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3927_ _1368_ _1590_ _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input297_I ic0_mem_data[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6646_ _0219_ clknet_leaf_24_core_clock dmmu0.page_table\[15\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3858_ immu_0.page_table\[0\]\[4\] immu_0.page_table\[1\]\[4\] immu_0.page_table\[2\]\[4\]
+ immu_0.page_table\[3\]\[4\] _1463_ _1391_ _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_41_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3229__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5543__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3789_ immu_0.page_table\[8\]\[2\] immu_0.page_table\[9\]\[2\] immu_0.page_table\[10\]\[2\]
+ immu_0.page_table\[11\]\[2\] _1424_ _1455_ _1457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6577_ _0150_ clknet_leaf_17_core_clock immu_0.page_table\[4\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_31_core_clock clknet_3_3_0_core_clock clknet_leaf_31_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5528_ _2645_ _0292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input60_I c0_o_req_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6099__A2 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5459_ immu_1.high_addr_off\[3\] _1852_ _2603_ _2607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput550 net550 dcache_mem_i_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput561 net561 dcache_mem_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput572 net572 dcache_wb_i_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput583 net583 ic0_mem_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_61_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3857__A1 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput594 net594 ic0_mem_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3857__B2 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7129_ net74 net597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5059__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_106_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6544__CLK clknet_leaf_18_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6023__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4034__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3468__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_2114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output683_I net683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_70_core_clock clknet_3_4_0_core_clock clknet_leaf_70_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7148__I net403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6694__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_56_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4273__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3076__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4830_ _2228_ _0011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4761_ _1817_ _2175_ _2177_ immu_0.page_table\[14\]\[8\] _2186_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_51_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3712_ _1381_ _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
X_6500_ _0073_ clknet_leaf_13_core_clock dmmu0.page_table\[14\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4692_ _2059_ _2139_ _2142_ net825 _2145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6431_ _0004_ clknet_leaf_108_core_clock immu_0.page_table\[13\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3643_ _1302_ net363 _1325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5525__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6362_ _0744_ clknet_leaf_75_core_clock immu_1.page_table\[12\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3574_ _1287_ net420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5313_ _2455_ _2516_ _2518_ dmmu0.page_table\[12\]\[3\] _2522_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6417__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6293_ _0675_ clknet_leaf_80_core_clock immu_1.page_table\[1\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_1276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5289__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5828__A2 _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5244_ _2328_ _2470_ _2472_ immu_0.page_table\[2\]\[8\] _2481_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold18 immu_1.page_table\[14\]\[8\] net752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold29 dmmu1.page_table\[10\]\[6\] net763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5175_ _2437_ _0147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4126_ net659 _0815_ net564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__6567__CLK clknet_leaf_18_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _1368_ _1716_ _1717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input212_I dcache_mem_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6005__A2 _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4016__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _2310_ _0058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4319__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6629_ _0202_ clknet_leaf_30_core_clock dmmu0.page_table\[12\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_2006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output431_I net431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3550__I0 net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3180__B _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4255__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4558__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3355__B _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4730__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3290_ _0882_ dmmu0.page_table\[12\]\[4\] _1036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_72_2373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3297__A2 _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3049__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6980_ _0553_ clknet_leaf_80_core_clock immu_1.page_table\[8\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4246__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ _2788_ _2873_ _2875_ dmmu1.page_table\[6\]\[4\] _2880_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_2177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5862_ _2782_ _2836_ _2838_ net833 _2840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4813_ _2217_ _0005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4549__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5746__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5793_ _2799_ _0403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4744_ _2176_ _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3852__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4675_ _2133_ _0760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6414_ _0796_ clknet_leaf_105_core_clock immu_0.page_table\[14\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3626_ _1316_ net698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3265__B _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3557_ _1278_ net549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6345_ _0727_ clknet_leaf_76_core_clock immu_1.page_table\[14\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input162_I c1_o_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6276_ _0658_ clknet_leaf_85_core_clock immu_1.page_table\[6\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3488_ _0875_ _1224_ _1226_ _0878_ _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_55_1870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput108 c1_o_c_instr_page net108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5227_ _2471_ _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput119 c1_o_mem_addr[10] net119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4485__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5682__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5158_ _2426_ _0141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_32_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input23_I c0_o_mem_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4109_ _1535_ net255 _1764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4237__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5089_ _2267_ _2382_ _2384_ immu_0.page_table\[7\]\[2\] _2387_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5434__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5985__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4788__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_1674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_1685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4115__I _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3212__A2 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output479_I net479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4960__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6732__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4173__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7161__I net175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6882__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3523__I0 _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_80_2631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_2030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_2041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5728__A1 _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ _2003_ _0675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_74_2424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6153__A1 _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold307 dmmu1.page_table\[12\]\[12\] net1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_46_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_2435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold318 dmmu0.page_table\[10\]\[3\] net1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3411_ _1149_ _1151_ _0878_ _1152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xhold329 dmmu0.page_table\[10\]\[7\] net1063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_68_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4391_ _1824_ _1957_ _1959_ net927 _1960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6130_ net559 _0818_ _2991_ _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_21_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3342_ dmmu1.page_table\[4\]\[7\] dmmu1.page_table\[5\]\[7\] dmmu1.page_table\[6\]\[7\]
+ dmmu1.page_table\[7\]\[7\] _0898_ _0909_ _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6061_ _2849_ _2941_ _2943_ net916 _2953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3273_ _0865_ dmmu0.page_table\[4\]\[4\] _1019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4467__A1 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4011__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5012_ _2342_ _0079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_1743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_2239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3690__A2 net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6963_ _0536_ clknet_leaf_54_core_clock dmmu1.page_table\[0\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5967__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_2038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5914_ _2869_ _0454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6605__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6894_ _0467_ clknet_leaf_66_core_clock dmmu1.page_table\[6\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5845_ _2829_ _0425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4078__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5776_ _2789_ _0396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_40_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6755__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4727_ _2165_ _0780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4942__A2 _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input377_I ic1_wb_adr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4658_ _1912_ _2122_ _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_57_1910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput90 c0_sr_bus_addr[8] net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3609_ _1303_ _1305_ _1307_ net703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_57_1932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4589_ _2065_ _2075_ _2077_ net853 _2083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_3_7_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_2047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6328_ _0710_ clknet_leaf_62_core_clock immu_1.page_table\[15\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_1807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6259_ _0641_ clknet_leaf_88_core_clock immu_1.page_table\[4\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3681__A2 net253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6285__CLK clknet_leaf_36_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4630__A1 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Right_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output596_I net596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5186__A2 _2429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4933__A2 _2285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7156__I net164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_20_Right_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5110__A2 _2397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6628__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5949__A1 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_2103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3960_ immu_1.page_table\[8\]\[7\] immu_1.page_table\[9\]\[7\] immu_1.page_table\[10\]\[7\]
+ immu_1.page_table\[11\]\[7\] _1441_ _1442_ _1623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_15_1624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6778__CLK clknet_leaf_99_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3891_ _1553_ _1554_ _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_2069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6171__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5630_ _1802_ _2699_ _2701_ dmmu0.page_table\[5\]\[3\] _2705_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3807__S0 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4924__A2 _2222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5561_ _2300_ _2663_ _2665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_60_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7066__I net406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4512_ _2034_ _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_48_1444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5492_ _2625_ _0276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold104 dmmu0.page_table\[11\]\[9\] net838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold115 dmmu1.page_table\[7\]\[7\] net849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold126 immu_0.page_table\[8\]\[9\] net860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4443_ _1819_ _1979_ _1982_ net874 _1992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold137 immu_1.page_table\[15\]\[0\] net871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_10_910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4688__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold148 immu_0.page_table\[4\]\[0\] net882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold159 immu_1.page_table\[9\]\[2\] net893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4374_ _1949_ _0643_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7162_ net176 net632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3325_ net150 dmmu1.long_off_reg\[0\] _1069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6113_ _1857_ _2975_ _2977_ dmmu1.page_table\[0\]\[5\] _2983_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7093_ net347 net500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3256_ _0899_ dmmu1.page_table\[8\]\[4\] _1002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6044_ _2944_ _0509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5101__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3112__A1 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3187_ dmmu0.page_table\[12\]\[1\] dmmu0.page_table\[13\]\[1\] dmmu0.page_table\[14\]\[1\]
+ dmmu0.page_table\[15\]\[1\] _0872_ _0868_ _0936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3663__A2 net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4860__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input125_I c1_o_mem_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _0519_ clknet_leaf_63_core_clock dmmu1.page_table\[2\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_27_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6877_ _0450_ clknet_leaf_54_core_clock dmmu1.page_table\[7\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_14_Left_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5168__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5828_ _2682_ _2818_ _2820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_14_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input90_I c0_sr_bus_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3179__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5759_ _2031_ _2137_ _2777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4915__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6117__A1 _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5340__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3351__A1 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold1_I ic0_wb_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5628__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output511_I net511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3654__A2 net247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4603__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5800__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_2009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5159__A2 _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4367__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6300__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_2097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6450__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3110_ net53 _0859_ _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_78_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ net117 immu_1.high_addr_off\[7\] _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5095__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3041_ net559 _0818_ _0819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3645__A2 net309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput280 ic0_mem_data[12] net280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput291 ic0_mem_data[22] net291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_1101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_63_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6800_ _0373_ clknet_leaf_41_core_clock dmmu1.page_table\[12\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4992_ _2329_ _0072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6731_ _0304_ clknet_leaf_96_core_clock dmmu0.page_table\[3\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3943_ _1606_ _1549_ _1607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6662_ _0235_ clknet_leaf_12_core_clock dmmu0.page_table\[11\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3874_ _1537_ _1538_ _1416_ _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_1498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _2694_ _0328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6593_ _0166_ clknet_leaf_5_core_clock immu_0.page_table\[2\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3257__C _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5544_ _2655_ _0298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_21_core_clock clknet_3_2_0_core_clock clknet_leaf_21_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3581__A1 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5475_ _2451_ _2613_ _2615_ dmmu0.page_table\[4\]\[1\] _2617_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_2115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4426_ _1983_ _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3333__A1 net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7145_ net400 net615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4357_ _1868_ _1927_ _1929_ immu_1.page_table\[5\]\[9\] _1939_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input242_I dcache_wb_adr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3308_ dmmu0.page_table\[12\]\[5\] dmmu0.page_table\[13\]\[5\] dmmu0.page_table\[14\]\[5\]
+ dmmu0.page_table\[15\]\[5\] _0872_ _0868_ _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7076_ net360 net513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4288_ _1899_ _0607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6943__CLK clknet_leaf_57_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3239_ dmmu1.page_table\[8\]\[3\] dmmu1.page_table\[9\]\[3\] dmmu1.page_table\[10\]\[3\]
+ dmmu1.page_table\[11\]\[3\] _0889_ _0931_ _0986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_39_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6027_ _2794_ _2924_ _2926_ net839 _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_2082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4833__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4597__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6929_ _0502_ clknet_leaf_56_core_clock dmmu1.page_table\[3\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_60_core_clock clknet_3_7_0_core_clock clknet_leaf_60_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4349__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__A2 _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output559_I net559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6473__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5313__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4521__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3911__B _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3627__A2 net270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3202__I _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3486__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5001__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3238__S1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6816__CLK clknet_leaf_40_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3590_ _1295_ net413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3563__A1 _1154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5260_ _2491_ _0178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3315__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6966__CLK clknet_leaf_57_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4211_ net201 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_76_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5191_ _2446_ _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_62_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4142_ net105 _1786_ _1787_ _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_4073_ immu_1.page_table\[4\]\[10\] immu_1.page_table\[5\]\[10\] immu_1.page_table\[6\]\[10\]
+ immu_1.page_table\[7\]\[10\] _1435_ _1469_ _1733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_21_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3174__S0 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6017__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4291__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6346__CLK clknet_leaf_75_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4579__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4975_ _2320_ _0064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5240__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6714_ _0287_ clknet_leaf_30_core_clock dmmu0.page_table\[13\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3926_ immu_0.page_table\[8\]\[6\] immu_0.page_table\[9\]\[6\] immu_0.page_table\[10\]\[6\]
+ immu_0.page_table\[11\]\[6\] _1424_ _1371_ _1590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_50_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6645_ _0218_ clknet_leaf_26_core_clock dmmu0.page_table\[15\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3857_ _1408_ _1521_ _1522_ net107 _1301_ _1523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_73_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3229__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input192_I c1_sr_bus_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5543__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6576_ _0149_ clknet_leaf_20_core_clock immu_0.page_table\[4\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3788_ immu_0.page_table\[0\]\[2\] immu_0.page_table\[1\]\[2\] immu_0.page_table\[2\]\[2\]
+ immu_0.page_table\[3\]\[2\] _1424_ _1455_ _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_6_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4751__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5527_ net95 _2629_ _2631_ dmmu0.page_table\[13\]\[12\] _2645_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6099__A3 _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput540 net540 dcache_mem_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5458_ _2606_ _0261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input53_I c0_o_mem_long_mode vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput551 net551 dcache_mem_i_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3306__A1 net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput562 net562 dcache_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput573 net573 dcache_wb_i_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4409_ _1868_ _1957_ _1959_ net755 _1969_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput584 net584 ic0_mem_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput595 net595 ic0_mem_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5389_ _2565_ _0233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3857__A2 _1521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7128_ net73 net596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5059__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3731__B _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7059_ net296 net447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5502__I _2631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4034__A2 _1694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3468__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6839__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3093__I0 net129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6989__CLK clknet_leaf_72_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3906__B _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7164__I net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6219__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6369__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4273__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4760_ _2185_ _0793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3711_ net385 _1380_ net2 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__3784__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ _2144_ _0765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6430_ _0003_ clknet_leaf_106_core_clock immu_0.page_table\[13\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3642_ _1324_ net691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5525__A2 _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6361_ _0743_ clknet_leaf_61_core_clock immu_1.page_table\[12\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7074__I net358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3573_ net223 _1204_ _1287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_49_Right_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_1233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5312_ _2521_ _0200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6292_ _0674_ clknet_leaf_82_core_clock immu_1.page_table\[1\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5289__A1 _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5243_ _2480_ _0172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold19 dmmu0.page_table\[6\]\[12\] net753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_23_1575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5174_ _2271_ _2430_ _2432_ net786 _2437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4125_ _1774_ net483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4056_ immu_0.page_table\[0\]\[10\] immu_0.page_table\[1\]\[10\] immu_0.page_table\[2\]\[10\]
+ immu_0.page_table\[3\]\[10\] _1370_ _1391_ _1716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_56_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_58_Right_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input205_I c1_sr_bus_data_o[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3777__I _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4016__A2 _1672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4958_ _2277_ _2299_ _2302_ dmmu0.page_table\[7\]\[7\] _2310_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3775__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3909_ _1377_ _1573_ _1574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_19_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4889_ _2262_ _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_69_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_43_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6628_ _0201_ clknet_leaf_26_core_clock dmmu0.page_table\[12\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Right_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4724__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6559_ _0132_ clknet_leaf_4_core_clock immu_0.page_table\[5\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6511__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3550__I1 net32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_76_Right_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4255__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6661__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7159__I net173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3310__S0 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5507__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_2_Left_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4191__A1 net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_2363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6191__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_1914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5930_ _2879_ _0460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_2178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5861_ _2839_ _0431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4812_ _1812_ _2208_ _2210_ net1047 _2217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5792_ _2047_ _2777_ _2779_ net750 _2799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5746__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4954__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4743_ _2140_ _2174_ _2176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4674_ _2069_ _2123_ _2125_ net762 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3509__A1 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6413_ _0795_ clknet_leaf_107_core_clock immu_0.page_table\[14\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4706__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3625_ _1308_ net269 _1316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6344_ _0726_ clknet_leaf_71_core_clock immu_1.page_table\[14\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3556_ net140 net35 _0841_ _1278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6534__CLK clknet_leaf_2_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6275_ _0657_ clknet_leaf_84_core_clock immu_1.page_table\[6\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3487_ _0877_ _1225_ _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_55_1860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input155_I c1_o_mem_high_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput109 c1_o_icache_flush net109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5226_ _1980_ _2469_ _2471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3368__S0 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4485__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5682__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6684__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5157_ _2330_ _2414_ _2416_ immu_0.page_table\[5\]\[9\] _2426_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_32_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input322_I ic0_wb_adr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4108_ _1761_ _1762_ _1763_ net702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_32_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5088_ _2386_ _0111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input16_I c0_o_mem_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4237__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5434__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4039_ net10 immu_0.high_addr_off\[5\] _1699_ _1700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_75_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3501__S _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5985__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_2044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3748__A1 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_2077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4131__I _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4173__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5370__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3920__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5122__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3987__A1 net113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_68_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6407__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_2031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3210__I net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__A2 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_2550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6557__CLK clknet_leaf_3_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_2414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6153__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_2425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold308 dmmu1.page_table\[4\]\[2\] net1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_29_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_2436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold319 immu_0.page_table\[2\]\[9\] net1053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3410_ _0877_ _1150_ _1151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3211__I0 _0956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ _1958_ _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_0_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3341_ dmmu1.page_table\[0\]\[7\] dmmu1.page_table\[1\]\[7\] dmmu1.page_table\[2\]\[7\]
+ dmmu1.page_table\[3\]\[7\] _0898_ _0901_ _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3813__C _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6060_ _2952_ _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3272_ dmmu0.page_table\[5\]\[4\] _1018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4467__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input8_I c0_o_instr_long_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4011__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5011_ _2267_ _2337_ _2339_ net947 _2342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_2011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6962_ _0535_ clknet_leaf_56_core_clock dmmu1.page_table\[0\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5967__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_2006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3978__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5913_ _2851_ _2855_ _2857_ dmmu1.page_table\[7\]\[10\] _2869_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6893_ _0466_ clknet_leaf_60_core_clock dmmu1.page_table\[6\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4216__I _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ _1814_ _2819_ _2821_ dmmu0.page_table\[1\]\[7\] _2829_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4078__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4927__B1 _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5775_ _2788_ _2778_ _2780_ dmmu1.page_table\[10\]\[4\] _2789_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_40_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4726_ _1809_ _2157_ _2159_ immu_0.page_table\[15\]\[5\] _2165_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_1073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4657_ _2122_ _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_70_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input272_I dcache_wb_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3608_ _1306_ net274 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput80 c0_sr_bus_addr[13] net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5352__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput91 c0_sr_bus_addr[9] net91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4588_ _2082_ _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3902__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6327_ _0709_ clknet_leaf_61_core_clock immu_1.page_table\[15\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3539_ _1269_ net555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3723__C _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6258_ _0640_ clknet_leaf_84_core_clock immu_1.page_table\[4\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5209_ _2459_ _2447_ _2449_ immu_0.page_table\[3\]\[5\] _2460_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_4_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6189_ _1796_ _3026_ _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3969__A1 net8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3513__S0 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4630__A2 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output491_I net491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_2084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3186__B _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7172__I net109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3406__S _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5646__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5949__A2 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3504__S0 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3890_ _1553_ _1554_ _1555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_2_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3875__I _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3807__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4385__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5560_ _2663_ _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_53_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4511_ _1980_ _2032_ _2034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_11_core_clock clknet_3_1_0_core_clock clknet_leaf_11_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5491_ _2529_ _2613_ _2615_ dmmu0.page_table\[4\]\[9\] _2625_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold105 dmmu1.page_table\[3\]\[7\] net839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold116 immu_1.page_table\[7\]\[4\] net850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4442_ _1991_ _0669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold127 immu_1.page_table\[12\]\[1\] net861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold138 dmmu1.page_table\[1\]\[7\] net872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold149 dmmu0.page_table\[9\]\[12\] net883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4688__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5885__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7161_ net175 net631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4373_ _1855_ _1942_ _1944_ net1026 _1949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_1191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6112_ _2982_ _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3324_ _1064_ _1065_ _1066_ _1067_ _0906_ _0912_ _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_7092_ net346 net499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6043_ _2776_ _2941_ _2943_ net747 _2944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3255_ dmmu1.page_table\[9\]\[4\] _1001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__3115__I _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3743__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3186_ _0931_ _0934_ _0884_ _0935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4860__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input118_I c1_o_mem_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _0518_ clknet_leaf_62_core_clock dmmu1.page_table\[2\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6722__CLK clknet_leaf_36_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5660__I1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_50_core_clock clknet_3_7_0_core_clock clknet_leaf_50_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_27_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6876_ _0449_ clknet_leaf_54_core_clock dmmu1.page_table\[7\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_27_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5827_ _2818_ _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_17_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5412__I1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3179__A2 _0927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6872__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ _1823_ _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5573__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input83_I c0_sr_bus_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4709_ _2153_ _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6117__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5689_ _2737_ _0361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4128__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_2090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3226__S _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3351__A2 net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5628__A1 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6252__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output504_I net504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__A2 _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6053__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5800__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_1295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4367__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5095__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3040_ mem_dcache_arb.req1_pending net159 _0809_ _0817_ _0818_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6745__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput270 dcache_wb_o_dat[8] net270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput281 ic0_mem_data[13] net281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput292 ic0_mem_data[23] net292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4991_ _2328_ _2317_ _2319_ dmmu0.page_table\[14\]\[8\] _2329_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_19_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6730_ _0303_ clknet_leaf_96_core_clock dmmu0.page_table\[3\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3942_ net111 immu_1.high_addr_off\[1\] _1606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6895__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6661_ _0234_ clknet_leaf_9_core_clock dmmu0.page_table\[11\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3873_ immu_1.page_table\[4\]\[5\] immu_1.page_table\[5\]\[5\] immu_1.page_table\[6\]\[5\]
+ immu_1.page_table\[7\]\[5\] _1435_ _1469_ _1538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_6_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7077__I net361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5612_ _2529_ _2681_ _2684_ net875 _2694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6592_ _0165_ clknet_leaf_4_core_clock immu_0.page_table\[2\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5543_ _2459_ _2647_ _2649_ net888 _2655_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5307__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3581__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5474_ _2616_ _0267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput700 net700 inner_wb_o_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_48_1286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5858__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4425_ _1777_ _1979_ _1982_ net766 _1983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6275__CLK clknet_leaf_84_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7144_ net399 net614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4356_ _1938_ _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3307_ _0934_ _1049_ _1050_ _1051_ _0841_ _1052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7075_ net359 net512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4287_ _1845_ _1894_ _1897_ immu_1.page_table\[0\]\[1\] _1899_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input235_I dcache_wb_adr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6026_ _2933_ _0502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3238_ dmmu1.page_table\[12\]\[3\] dmmu1.page_table\[13\]\[3\] dmmu1.page_table\[14\]\[3\]
+ dmmu1.page_table\[15\]\[3\] _0889_ _0931_ _0985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4833__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3169_ _0907_ _0918_ _0919_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input402_I inner_wb_i_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6035__A1 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4597__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6928_ _0501_ clknet_leaf_55_core_clock dmmu1.page_table\[3\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6859_ _0432_ clknet_leaf_48_core_clock dmmu1.page_table\[8\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4349__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6618__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output454_I net454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4521__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3955__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4521__B2 dmmu1.page_table\[14\]\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6768__CLK clknet_leaf_40_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output621_I net621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3911__C _1575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3260__A1 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5537__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5001__A2 _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_2097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6298__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3563__A2 _1186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4210_ _1844_ _0584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3166__I2 dmmu1.page_table\[14\]\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _1789_ _2445_ _2446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_23_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4141_ net89 net88 net87 _1787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__6177__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4072_ net107 _1730_ _1731_ _1732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_56_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3174__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6017__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4579__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4974_ _2258_ _2317_ _2319_ dmmu0.page_table\[14\]\[0\] _2320_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_1_core_clock clknet_3_0_0_core_clock clknet_leaf_1_core_clock vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5240__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3925_ _1375_ _1588_ _1589_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6713_ _0286_ clknet_leaf_34_core_clock dmmu0.page_table\[13\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3251__A1 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_108_core_clock clknet_3_0_0_core_clock clknet_leaf_108_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__I _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6644_ _0217_ clknet_leaf_35_core_clock dmmu0.page_table\[15\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3856_ net110 immu_1.high_addr_off\[0\] _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6575_ _0148_ clknet_leaf_20_core_clock immu_0.page_table\[4\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3787_ net313 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_60_1995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4751__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input185_I c1_sr_bus_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5526_ _2644_ _0291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6910__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5457_ immu_1.high_addr_off\[2\] _1849_ _2603_ _2606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput530 net530 dcache_mem_addr[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput541 net541 dcache_mem_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput552 net552 dcache_mem_i_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input352_I ic1_mem_data[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput563 net563 dcache_rst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4408_ _1968_ _0658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4503__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput574 net574 dcache_wb_i_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_22_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5388_ _2529_ _2553_ _2555_ net838 _2565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput585 net585 ic0_mem_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_61_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input46_I c0_o_mem_high_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput596 net596 ic0_mem_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7127_ net72 net595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4339_ _1824_ _1927_ _1929_ immu_1.page_table\[5\]\[0\] _1930_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5059__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7058_ net295 net446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3731__C _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4267__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6009_ _1874_ _1891_ _2030_ _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_55_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3242__A1 _0974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3093__I1 net24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6440__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7180__I net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3710_ net3 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_51_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3784__A2 _1427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4690_ _2057_ _2139_ _2142_ immu_1.page_table\[10\]\[1\] _2144_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_0_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3641_ _0812_ net262 _1324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_43_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_2093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6360_ _0742_ clknet_leaf_61_core_clock immu_1.page_table\[12\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3572_ _1286_ net419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5311_ _2453_ _2516_ _2518_ net816 _2521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_1977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6291_ _0673_ clknet_leaf_98_core_clock dmmu0.page_table\[0\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_75_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5289__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3919__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5242_ _2463_ _2470_ _2472_ net1010 _2480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4497__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5173_ _2436_ _0146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4124_ net213 _0831_ _1774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6313__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 c0_o_c_data_page net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_78_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4055_ _1375_ _1714_ _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3847__I0 net237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5997__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3472__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6463__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input100_I c0_sr_bus_data_o[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ _2309_ _0057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3908_ _1563_ _1566_ _1569_ _1572_ _1573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3775__A2 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4972__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4888_ _1980_ _2260_ _2262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_7_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6627_ _0200_ clknet_leaf_26_core_clock dmmu0.page_table\[12\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3839_ immu_1.page_table\[12\]\[3\] immu_1.page_table\[13\]\[3\] _1474_ _1506_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4724__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ _0131_ clknet_leaf_7_core_clock immu_0.page_table\[6\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5509_ _2455_ _2630_ _2632_ net866 _2636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6489_ _0062_ clknet_leaf_11_core_clock dmmu0.page_table\[7\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4660__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6956__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3310__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7175__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6336__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6486__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_2179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5860_ _2776_ _2836_ _2838_ net957 _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4811_ _2216_ _0004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_2079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5791_ _2798_ _0402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4403__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4954__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4742_ _2174_ _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_7_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4673_ _2132_ _0759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6412_ _0794_ clknet_leaf_107_core_clock immu_0.page_table\[14\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3624_ _1315_ net697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4706__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5903__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6343_ _0725_ clknet_leaf_74_core_clock immu_1.page_table\[14\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3555_ _1277_ net548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3118__I _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6274_ _0656_ clknet_leaf_87_core_clock immu_1.page_table\[6\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3486_ dmmu0.page_table\[0\]\[11\] dmmu0.page_table\[1\]\[11\] dmmu0.page_table\[2\]\[11\]
+ dmmu0.page_table\[3\]\[11\] _0871_ _0866_ _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_55_1850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5225_ _2469_ _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_55_1861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3368__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6829__CLK clknet_leaf_68_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input148_I c1_o_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5682__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5156_ _2425_ _0140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_51_1747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3693__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4890__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4107_ _1535_ net273 _1763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5087_ _2265_ _2382_ _2384_ immu_0.page_table\[7\]\[1\] _2386_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_32_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input315_I ic0_wb_adr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5434__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4038_ _1666_ _1697_ _1698_ _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6979__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4642__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_1676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5989_ _2786_ _2907_ _2909_ net910 _2913_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3748__A2 _1417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6147__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5370__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4173__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3920__A2 _1583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3684__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3698__I _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_2633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_2032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_2562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_2415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_2426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold309 dmmu1.page_table\[13\]\[12\] net1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_74_2437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3340_ net152 dmmu1.long_off_reg\[2\] _1082_ _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_61_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3271_ dmmu0.page_table\[6\]\[4\] dmmu0.page_table\[7\]\[4\] _0872_ _1017_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5010_ _2341_ _0078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4872__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6185__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6961_ _0534_ clknet_leaf_62_core_clock dmmu1.page_table\[1\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3427__A1 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5912_ _2868_ _0453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_40_core_clock clknet_3_6_0_core_clock clknet_leaf_40_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6892_ _0465_ clknet_leaf_58_core_clock dmmu1.page_table\[6\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ _2828_ _0424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4927__A1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4927__B2 _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5774_ _1854_ _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_40_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6501__CLK clknet_leaf_10_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4725_ _2164_ _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4232__I _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4656_ _1826_ _1839_ _1874_ _2122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_47_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput70 c0_o_req_addr[5] net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3607_ inner_wb_arbiter.o_sel_sig _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_47_1159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput81 c0_sr_bus_addr[14] net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5352__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4587_ _2063_ _2075_ _2077_ immu_1.page_table\[14\]\[4\] _2082_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_57_1923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput92 c0_sr_bus_data_o[0] net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6651__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input265_I dcache_wb_o_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3538_ net146 net41 _1267_ _1269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6326_ _0708_ clknet_leaf_68_core_clock dmmu1.page_table\[14\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3292__B _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6257_ _0639_ clknet_leaf_82_core_clock immu_1.page_table\[4\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3469_ _0907_ _1207_ _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5208_ _1808_ _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_42_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6188_ _1781_ _1788_ _2284_ _3026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_4_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3666__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5139_ _2258_ _2414_ _2416_ immu_0.page_table\[5\]\[0\] _2417_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3418__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4615__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3513__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4630__A3 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output484_I net484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Left_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5646__A2 _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3657__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3930__B _1593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_2230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Left_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5949__A3 _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6071__A2 _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3504__S1 net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4082__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6524__CLK clknet_leaf_2_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4510_ _2032_ _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_53_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6674__CLK clknet_leaf_36_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5490_ _2624_ _0275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Left_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_14_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5334__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold106 dmmu1.page_table\[6\]\[11\] net840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4441_ _1817_ _1979_ _1982_ dmmu0.page_table\[0\]\[8\] _1991_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold117 dmmu0.page_table\[6\]\[1\] net851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_9_Right_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold128 dmmu1.page_table\[11\]\[11\] net862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_10_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold139 dmmu1.page_table\[9\]\[7\] net873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7160_ net174 net630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4372_ _1948_ _0642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3896__A1 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6111_ _1854_ _2975_ _2977_ dmmu1.page_table\[0\]\[4\] _2982_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3323_ dmmu1.page_table\[8\]\[6\] dmmu1.page_table\[9\]\[6\] dmmu1.page_table\[10\]\[6\]
+ dmmu1.page_table\[11\]\[6\] _0888_ _0901_ _1067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7091_ net345 net498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6042_ _2942_ _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3254_ dmmu1.page_table\[10\]\[4\] dmmu1.page_table\[11\]\[4\] _0908_ _1000_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3648__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4936__B _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4845__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3743__S1 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3185_ net124 _0932_ _0892_ _0933_ _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_59_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_53_Left_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_1731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6944_ _0517_ clknet_leaf_58_core_clock dmmu1.page_table\[2\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6875_ _0448_ clknet_leaf_65_core_clock dmmu1.page_table\[7\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5826_ _1976_ _2484_ _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_14_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3287__B _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5573__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ _2775_ _0391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input382_I ic1_wb_stb vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_62_Left_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4708_ _2105_ _2138_ _2141_ immu_1.page_table\[10\]\[10\] _2153_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5688_ _2101_ _2726_ _2728_ dmmu1.page_table\[13\]\[8\] _2737_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input76_I c0_sr_bus_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4128__A2 net230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4639_ _2113_ _0744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3887__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3431__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6309_ _0691_ clknet_leaf_80_core_clock immu_1.page_table\[3\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5089__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5628__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3639__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_71_Left_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6547__CLK clknet_leaf_8_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6053__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4064__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5261__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5800__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3811__A1 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_3_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5013__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Left_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3197__B _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4367__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_5_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7183__I net402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3422__S0 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_2107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput260 dcache_wb_o_dat[13] net260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput271 dcache_wb_o_dat[9] net271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput282 ic0_mem_data[14] net282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput293 ic0_mem_data[24] net293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4055__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4990_ net103 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3102__I0 net133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3941_ _1408_ _1599_ _1604_ _1605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_50_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3872_ immu_1.page_table\[0\]\[5\] immu_1.page_table\[1\]\[5\] immu_1.page_table\[2\]\[5\]
+ immu_1.page_table\[3\]\[5\] _1435_ _1469_ _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6660_ _0233_ clknet_leaf_12_core_clock dmmu0.page_table\[11\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5611_ _2693_ _0327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5555__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6591_ _0164_ clknet_leaf_10_core_clock immu_0.page_table\[3\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5542_ _2654_ _0297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5307__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ _2444_ _2613_ _2615_ dmmu0.page_table\[4\]\[0\] _2616_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput701 net701 inner_wb_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4510__I _2032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3318__B1 _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4424_ _1981_ _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_26_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4355_ _1866_ _1927_ _1929_ net791 _1938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7143_ net398 net613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3126__I _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3306_ net158 _0893_ _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7074_ net358 net511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4286_ _1890_ _1894_ _1897_ _1898_ _0606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4818__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3237_ _0982_ _0983_ _0842_ _0984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6025_ _2792_ _2924_ _2926_ dmmu1.page_table\[3\]\[6\] _2933_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input130_I c1_o_mem_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5491__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input228_I dcache_mem_o_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3168_ dmmu1.page_table\[8\]\[0\] dmmu1.page_table\[9\]\[0\] dmmu1.page_table\[10\]\[0\]
+ dmmu1.page_table\[11\]\[0\] _0899_ _0902_ _0918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_74_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6035__A2 _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3099_ _0852_ net539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4046__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_82_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4597__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5794__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6927_ _0500_ clknet_leaf_56_core_clock dmmu1.page_table\[3\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3729__C _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6858_ _0431_ clknet_leaf_47_core_clock dmmu1.page_table\[8\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_1955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5809_ _2809_ _0409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4349__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6789_ _0362_ clknet_leaf_66_core_clock dmmu1.page_table\[13\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3404__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output447_I net447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4521__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3955__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_2015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4037__A1 net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5234__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7178__I net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3260__A2 dmmu1.page_table\[14\]\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_2019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3563__A3 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6712__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4140_ net86 _1786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4071_ _1726_ _1729_ _1731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6862__CLK clknet_leaf_48_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5473__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6017__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4973_ _2318_ _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_1387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6712_ _0285_ clknet_leaf_25_core_clock dmmu0.page_table\[13\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3924_ immu_0.page_table\[12\]\[6\] immu_0.page_table\[13\]\[6\] immu_0.page_table\[14\]\[6\]
+ immu_0.page_table\[15\]\[6\] _1424_ _1455_ _1588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_46_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6643_ _0216_ clknet_leaf_25_core_clock dmmu0.page_table\[15\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3855_ _1517_ _1520_ _1440_ _1521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6242__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3786_ _1454_ net664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6574_ _0147_ clknet_leaf_18_core_clock immu_0.page_table\[4\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_60_1996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5525_ net94 _2629_ _2631_ net806 _2644_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4751__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input178_I c1_o_req_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3284__C _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput520 net520 dcache_mem_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_14_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5456_ _2605_ _0260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6392__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput531 net531 dcache_mem_addr[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput542 net542 dcache_mem_cache_enable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput553 net553 dcache_mem_i_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4407_ _1866_ _1957_ _1959_ net1009 _1968_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput564 net564 dcache_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__5700__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput575 net575 dcache_wb_i_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5387_ _2564_ _0232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput586 net586 ic0_mem_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_61_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input345_I ic1_mem_data[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7126_ net71 net594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput597 net597 ic0_mem_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4338_ _1928_ _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input39_I c0_o_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7057_ net294 net445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4269_ _1864_ _1876_ _1878_ immu_1.page_table\[7\]\[7\] _1886_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4267__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6008_ _2922_ _0495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4019__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3242__A2 _0979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3873__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3475__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6735__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output564_I net564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6885__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6265__CLK clknet_leaf_84_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3864__S0 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3784__A3 _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3640_ _1323_ net690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3571_ net222 _1204_ _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5310_ _2520_ _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6290_ _0672_ clknet_leaf_98_core_clock dmmu0.page_table\[0\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5241_ _2479_ _0171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3919__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4497__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4041__S0 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3544__I0 net149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5172_ _2269_ _2430_ _2432_ net1039 _2436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4123_ _1773_ net466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_1599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 c0_o_c_instr_long net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4054_ immu_0.page_table\[4\]\[10\] immu_0.page_table\[5\]\[10\] immu_0.page_table\[6\]\[10\]
+ immu_0.page_table\[7\]\[10\] _1370_ _1391_ _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5997__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6608__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4235__I net207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3279__C _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4956_ _2275_ _2299_ _2302_ dmmu0.page_table\[7\]\[6\] _2309_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6758__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3907_ _1570_ _1571_ _1366_ _1572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4972__A2 _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4887_ _2260_ _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input295_I ic0_mem_data[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6626_ _0199_ clknet_leaf_25_core_clock dmmu0.page_table\[12\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3838_ _1440_ _1504_ _1505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6557_ _0130_ clknet_leaf_3_core_clock immu_0.page_table\[6\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5921__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3769_ _1437_ _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_70_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5508_ _2635_ _0282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6488_ _0061_ clknet_leaf_11_core_clock dmmu0.page_table\[7\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5439_ _2594_ _0254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3515__S _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7109_ net400 net577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6288__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4660__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output681_I net681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6165__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_2490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_19_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7191__I net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A1 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_2376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5676__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5428__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5979__A1 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_core_clock clknet_3_3_0_core_clock clknet_leaf_30_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_76_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6900__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4810_ _1809_ _2208_ _2210_ immu_0.page_table\[13\]\[5\] _2216_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4403__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5790_ _2105_ _2777_ _2779_ net765 _2798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5600__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3837__S0 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4741_ _1790_ _2173_ _2174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4954__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4672_ _2067_ _2123_ _2125_ net854 _2132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_12_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6411_ _0793_ clknet_leaf_106_core_clock immu_0.page_table\[14\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5903__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3623_ _1308_ net268 _1315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4706__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6342_ _0724_ clknet_leaf_76_core_clock immu_1.page_table\[14\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3554_ net139 net34 _1267_ _1277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6273_ _0655_ clknet_leaf_88_core_clock immu_1.page_table\[6\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3485_ dmmu0.page_table\[4\]\[11\] dmmu0.page_table\[5\]\[11\] dmmu0.page_table\[6\]\[11\]
+ dmmu0.page_table\[7\]\[11\] _0864_ _0867_ _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_11_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5224_ _1789_ _2468_ _2469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_55_1862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_1726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6430__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3134__I _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5155_ _2328_ _2414_ _2416_ net771 _2425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_51_1748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3693__A2 net311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4890__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4106_ _1350_ net327 _1360_ _1762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_32_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5086_ _2385_ _0110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4037_ net9 immu_0.high_addr_off\[4\] _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_21_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input210_I c1_sr_bus_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4642__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input308_I ic0_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6580__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_49_1677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5988_ _2912_ _0485_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4939_ _1977_ _2297_ _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_34_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6147__A1 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6609_ _0182_ clknet_leaf_16_core_clock immu_0.page_table\[1\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5370__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3220__I2 dmmu1.page_table\[14\]\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3381__A1 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5122__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3133__A1 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output527_I net527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3044__I _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3684__A2 net324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6923__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6083__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5830__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_2612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5189__A2 _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3819__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4397__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7186__I net390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6303__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4149__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_2416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5897__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_2427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_2438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3372__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6453__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3382__C _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3270_ _1014_ _0858_ _1015_ _1016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_20_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4321__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4872__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6960_ _0533_ clknet_leaf_64_core_clock dmmu1.page_table\[1\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5911_ _2849_ _2856_ _2858_ net787 _2868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6891_ _0464_ clknet_leaf_58_core_clock dmmu1.page_table\[6\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5842_ _1811_ _2819_ _2821_ dmmu0.page_table\[1\]\[6\] _2828_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_87_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5773_ _2787_ _0395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4927__A2 _2285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6129__A1 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4724_ _1806_ _2157_ _2159_ immu_0.page_table\[15\]\[4\] _2164_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_20_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4655_ _2121_ _0752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3129__I _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3606_ _0814_ net328 net659 _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput60 c0_o_req_addr[10] net60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput71 c0_o_req_addr[6] net71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5352__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput82 c0_sr_bus_addr[15] net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4586_ _2081_ _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_57_1924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput93 c0_sr_bus_data_o[10] net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_60_2039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6325_ _0707_ clknet_leaf_39_core_clock dmmu1.page_table\[14\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3537_ _1268_ net554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input160_I c1_o_mem_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input258_I dcache_wb_o_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6256_ _0638_ clknet_leaf_93_core_clock immu_1.page_table\[5\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3468_ dmmu1.page_table\[8\]\[11\] dmmu1.page_table\[9\]\[11\] dmmu1.page_table\[10\]\[11\]
+ dmmu1.page_table\[11\]\[11\] _0898_ _0901_ _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5207_ _2458_ _0158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6187_ net736 _3025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3399_ net48 dmmu0.long_off_reg\[3\] _1140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3666__A2 net320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5138_ _2415_ _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input21_I c0_o_mem_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ _2273_ _2367_ _2369_ immu_0.page_table\[8\]\[5\] _2375_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4615__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5812__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6326__CLK clknet_leaf_68_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4379__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5455__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6476__CLK clknet_leaf_102_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3106__A1 net50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4303__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3657__A2 net318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3930__C _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_2220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_2106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_2039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5031__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6819__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3593__A1 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4790__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4440_ _1990_ _0668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold107 immu_1.page_table\[4\]\[3\] net841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5334__A2 _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold118 immu_0.page_table\[4\]\[7\] net852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold129 immu_1.page_table\[10\]\[6\] net863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6969__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3345__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4371_ _1852_ _1942_ _1944_ net841 _1948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6110_ _2981_ _0538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3322_ dmmu1.page_table\[12\]\[6\] dmmu1.page_table\[13\]\[6\] dmmu1.page_table\[14\]\[6\]
+ dmmu1.page_table\[15\]\[6\] _0888_ _0901_ _1066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7090_ net344 net497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4001__C _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6041_ _1770_ _2940_ _2942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3253_ _0931_ _0995_ _0998_ _0896_ _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_20_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3648__A2 net370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4845__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3184_ net106 _0932_ _0933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__6047__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4508__I _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6943_ _0516_ clknet_leaf_57_core_clock dmmu1.page_table\[2\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6874_ _0447_ clknet_leaf_52_core_clock dmmu1.page_table\[7\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_27_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5825_ _2817_ _0417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6499__CLK clknet_leaf_21_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5756_ _2049_ _2759_ _2761_ dmmu1.page_table\[11\]\[12\] _2775_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5573__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4707_ _2152_ _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5687_ _2736_ _0360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input375_I ic1_wb_adr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4638_ _2059_ _2108_ _2110_ immu_1.page_table\[12\]\[2\] _2113_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input69_I c0_o_req_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4569_ _1866_ _2053_ _2055_ net931 _2071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3887__A2 _1546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3431__S1 _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6308_ _0690_ clknet_leaf_86_core_clock immu_1.page_table\[3\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5089__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6239_ _0621_ clknet_leaf_81_core_clock immu_1.page_table\[2\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3639__A2 net261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3523__S _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3195__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4064__A2 _1723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5261__A1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output594_I net594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5013__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3575__A1 net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4772__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3327__A1 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4102__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3422__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3433__S _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4827__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput250 dcache_wb_adr[5] net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput261 dcache_wb_o_dat[14] net261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6029__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput272 dcache_wb_sel[0] net272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput283 ic0_mem_data[15] net283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput294 ic0_mem_data[25] net294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3102__I1 net28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6641__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3940_ _1446_ _1601_ _1603_ _1604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_14_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3871_ _1306_ _1523_ _1534_ _1536_ net667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_58_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5610_ _2527_ _2681_ _2684_ net1028 _2693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5555__A2 _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6590_ _0163_ clknet_leaf_6_core_clock immu_0.page_table\[3\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6791__CLK clknet_leaf_40_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4763__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5541_ _2457_ _2647_ _2649_ dmmu0.page_table\[3\]\[4\] _2654_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5307__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5472_ _2614_ _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3318__A1 _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput702 net702 inner_wb_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4423_ _1980_ _1978_ _1981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4515__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3318__B2 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7142_ net397 net612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4354_ _1937_ _0635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_18_Left_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3305_ net150 dmmu1.long_off_reg\[0\] _1050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7073_ net357 net510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4285_ net737 _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3343__S _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4818__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ _2932_ _0501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3236_ _0915_ _0895_ _0983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_1903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_2074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5491__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3167_ _0897_ _0916_ _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input123_I c1_o_mem_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3098_ net131 net26 _0850_ _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4046__A2 net244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6926_ _0499_ clknet_leaf_51_core_clock dmmu1.page_table\[3\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _0430_ clknet_leaf_98_core_clock dmmu0.page_table\[1\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5808_ _2788_ _2802_ _2804_ dmmu1.page_table\[9\]\[4\] _2809_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6788_ _0361_ clknet_leaf_43_core_clock dmmu1.page_table\[13\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5739_ _2766_ _0382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_2018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3309__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3404__S1 _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6514__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3168__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_2038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6664__CLK clknet_leaf_104_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3052__I _0826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5234__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3096__I0 net130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3796__A1 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_2055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4745__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6194__CLK clknet_leaf_8_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5170__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4070_ _1726_ _1729_ _1730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5473__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3087__I0 net126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_26_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4972_ _2300_ _2316_ _2318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _0284_ clknet_leaf_30_core_clock dmmu0.page_table\[13\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3331__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4984__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3923_ _1383_ _1584_ _1586_ _1587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_54_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6642_ _0215_ clknet_leaf_29_core_clock dmmu0.page_table\[15\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3854_ _1518_ _1519_ _1446_ _1520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6573_ _0146_ clknet_leaf_20_core_clock immu_0.page_table\[4\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3785_ net235 _1453_ _1360_ _1454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5524_ _2643_ _0290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6537__CLK clknet_leaf_4_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ immu_1.high_addr_off\[1\] _1846_ _2603_ _2605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput510 net510 c1_i_req_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3137__I _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput521 net521 dcache_mem_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput532 net532 dcache_mem_addr[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput543 net543 dcache_mem_i_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_4406_ _1967_ _0657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput554 net554 dcache_mem_i_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_2095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5386_ _2527_ _2553_ _2555_ dmmu0.page_table\[11\]\[8\] _2564_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput565 net565 dcache_wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_41_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput576 net576 dcache_wb_i_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7125_ net70 net593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3711__A1 net385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput587 net587 ic0_mem_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4337_ _1912_ _1926_ _1928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput598 net598 ic0_mem_cache_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__6687__CLK clknet_leaf_91_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input240_I dcache_wb_adr[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input338_I ic1_mem_data[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7056_ net293 net444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_5_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4268_ _1885_ _0601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4267__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6007_ net200 _2906_ _2908_ dmmu1.page_table\[4\]\[12\] _2922_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3219_ dmmu1.page_table\[4\]\[2\] dmmu1.page_table\[5\]\[2\] dmmu1.page_table\[6\]\[2\]
+ dmmu1.page_table\[7\]\[2\] _0889_ _0931_ _0967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_39_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4199_ _1830_ net196 _1833_ _1834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_74_1635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4019__A2 net243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3600__I _1300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_2044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3778__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3322__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6909_ _0482_ clknet_leaf_63_core_clock dmmu1.page_table\[5\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3873__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3950__A1 net112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_2015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold290 dmmu0.page_table\[13\]\[8\] net1024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20_core_clock clknet_3_2_0_core_clock clknet_leaf_20_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_77_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7189__I net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3864__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3666__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4718__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4194__A1 _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3570_ _1285_ net418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3941__A1 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5240_ _2461_ _2470_ _2472_ immu_0.page_table\[2\]\[6\] _2479_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4497__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4041__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5694__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3544__I1 net44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Right_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5171_ _2435_ _0145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4122_ net212 _0831_ _1773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5446__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4249__A2 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4053_ _1708_ _1711_ _1579_ _1713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_21_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 c0_o_c_instr_page net3 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5997__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ _2308_ _0056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Right_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3906_ _1396_ immu_0.page_table\[9\]\[5\] _1390_ _1571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4886_ _1977_ _2259_ _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_74_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6625_ _0198_ clknet_leaf_25_core_clock dmmu0.page_table\[12\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3837_ immu_1.page_table\[8\]\[3\] immu_1.page_table\[9\]\[3\] immu_1.page_table\[10\]\[3\]
+ immu_1.page_table\[11\]\[3\] _1474_ _1469_ _1504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_34_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input190_I c1_sr_bus_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input288_I ic0_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6556_ _0129_ clknet_leaf_18_core_clock immu_0.page_table\[6\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5382__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3768_ _1434_ _1436_ net705 _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5921__A2 _2872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5507_ _2453_ _2630_ _2632_ net1083 _2635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3932__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6487_ _0060_ clknet_leaf_38_core_clock dmmu0.page_table\[7\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3699_ net312 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_63_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5438_ _2529_ _2582_ _2584_ net757 _2594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_36_Right_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input51_I c0_o_mem_high_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5369_ _2554_ _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7108_ net399 net576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_94_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7039_ net306 net457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3531__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3999__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4660__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Right_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4948__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6702__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6852__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3923__A1 _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Right_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_76_2480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_2491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A2 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5676__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5428__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6232__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5979__A2 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Right_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_2004 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6382__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5600__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3837__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4740_ _2154_ _2172_ _2173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_51_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ _2131_ _0758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6410_ _0792_ clknet_leaf_109_core_clock immu_0.page_table\[14\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3622_ _1314_ net696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_42_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_72_Right_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5903__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3914__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6341_ _0723_ clknet_leaf_71_core_clock immu_1.page_table\[14\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3553_ _1276_ net547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5116__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6272_ _0654_ clknet_leaf_84_core_clock immu_1.page_table\[6\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3843__C _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3484_ _0877_ _1220_ _1222_ _0958_ _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_42_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5223_ _1971_ _2172_ _2468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_55_1852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5154_ _2424_ _0139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_36_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4105_ _1348_ net381 _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4890__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5085_ _2258_ _2382_ _2384_ immu_0.page_table\[7\]\[0\] _2385_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4036_ net9 immu_0.high_addr_off\[4\] _1697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6725__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4642__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3150__I net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input203_I c1_sr_bus_data_o[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5987_ _2784_ _2907_ _2909_ net1042 _2912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6875__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4938_ _1780_ _2296_ _2297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_5_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input99_I c0_sr_bus_data_o[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6147__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4869_ _2250_ _0028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6608_ _0181_ clknet_leaf_17_core_clock immu_0.page_table\[1\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3905__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6539_ _0112_ clknet_leaf_3_core_clock immu_0.page_table\[7\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6255__CLK clknet_leaf_83_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6083__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3516__S0 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Left_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4156__I _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5830__A1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3060__I _0830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_2034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3819__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4397__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5594__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_2081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4149__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_2542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5346__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5897__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_2417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_74_2428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_2439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4321__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6748__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4872__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_1460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6898__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5910_ _2867_ _0452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6890_ _0463_ clknet_leaf_54_core_clock dmmu1.page_table\[6\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5841_ _2827_ _0423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_1477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5772_ _2786_ _2778_ _2780_ dmmu1.page_table\[10\]\[3\] _2787_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4723_ _2163_ _0778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_40_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6129__A2 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4654_ _2105_ _2107_ _2109_ immu_1.page_table\[12\]\[10\] _2121_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput50 c0_o_mem_high_addr[5] net50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3605_ _1304_ net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_47_1139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput61 c0_o_req_addr[11] net61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6278__CLK clknet_leaf_92_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput72 c0_o_req_addr[7] net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4585_ _2061_ _2075_ _2077_ immu_1.page_table\[14\]\[3\] _2081_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_57_1914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput83 c0_sr_bus_addr[1] net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_57_1925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput94 c0_sr_bus_data_o[11] net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6324_ _0706_ clknet_leaf_69_core_clock dmmu1.page_table\[14\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3994__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3536_ net145 net40 _1267_ _1268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6255_ _0637_ clknet_leaf_83_core_clock immu_1.page_table\[5\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3467_ _0897_ _1205_ _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_1762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input153_I c1_o_mem_high_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5206_ _2457_ _2447_ _2449_ immu_0.page_table\[3\]\[4\] _2458_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6186_ _3024_ _0571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3398_ _1118_ _1124_ _1139_ net528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_4_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5137_ _1980_ _2413_ _2415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3081__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input320_I ic0_wb_adr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6065__A1 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5068_ _2374_ _0103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5812__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input14_I c0_o_mem_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4615__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4019_ net659 net243 _1681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_2109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Right_0 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4379__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3051__A1 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4303__A1 net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3106__A2 net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_2210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5654__I1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_2107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3290__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5406__I1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__CLK clknet_leaf_108_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5319__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3593__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold108 dmmu0.page_table\[3\]\[0\] net842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold119 immu_1.page_table\[14\]\[5\] net853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4542__A1 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4370_ _1947_ _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6570__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3321_ dmmu1.page_table\[0\]\[6\] dmmu1.page_table\[1\]\[6\] dmmu1.page_table\[2\]\[6\]
+ dmmu1.page_table\[3\]\[6\] _0888_ _0910_ _1065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_10_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6040_ _2940_ _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3252_ _0889_ _0996_ _0997_ _0902_ _0998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_28_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I c0_o_instr_long_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4845__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3183_ net158 _0932_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__6047__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6942_ _0515_ clknet_leaf_56_core_clock dmmu1.page_table\[2\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6873_ _0446_ clknet_leaf_50_core_clock dmmu1.page_table\[7\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5824_ _2049_ _2801_ _2803_ net810 _2817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5755_ _2774_ _0390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4706_ _2103_ _2139_ _2142_ immu_1.page_table\[10\]\[9\] _2152_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5686_ _2069_ _2726_ _2728_ dmmu1.page_table\[13\]\[7\] _2736_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6913__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4637_ _2112_ _0743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input270_I dcache_wb_o_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4533__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3336__A2 _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input368_I ic1_wb_adr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4568_ _2070_ _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6307_ _0689_ clknet_leaf_79_core_clock immu_1.page_table\[3\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3519_ _0896_ _1256_ _1257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4499_ _1866_ _2014_ _2016_ immu_1.page_table\[3\]\[8\] _2025_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3804__S _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5089__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6238_ _0620_ clknet_leaf_91_core_clock immu_1.page_table\[2\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4297__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6169_ _2029_ _2601_ _3015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3195__S1 _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3895__I0 _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5261__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6443__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5549__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5013__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output587_I net587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4221__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3575__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6593__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3327__A2 _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3958__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4827__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput240 dcache_wb_adr[18] net240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput251 dcache_wb_adr[6] net251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6029__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput262 dcache_wb_o_dat[15] net262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput273 dcache_wb_sel[1] net273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput284 ic0_mem_data[16] net284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput295 ic0_mem_data[26] net295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5788__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3263__A1 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Left_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3870_ _1535_ net238 _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4763__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5540_ _2653_ _0296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5471_ _2300_ _2612_ _2614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_14_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput703 net703 inner_wb_stb vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4515__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4422_ _1769_ _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_48_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4515__B2 dmmu1.page_table\[14\]\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5712__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7141_ net396 net611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4353_ _1864_ _1927_ _1929_ net920 _1937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3304_ _0915_ _1042_ _1044_ _1046_ _1048_ _1049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_7072_ net356 net509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4284_ _1896_ _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6316__CLK clknet_leaf_69_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4818__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6023_ _2790_ _2924_ _2926_ net748 _2932_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3235_ _0980_ _0981_ _0907_ _0982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_1131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_99_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5491__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3166_ dmmu1.page_table\[12\]\[0\] dmmu1.page_table\[13\]\[0\] dmmu1.page_table\[14\]\[0\]
+ dmmu1.page_table\[15\]\[0\] _0899_ _0902_ _0916_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_78_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6466__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3097_ _0851_ net538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input116_I c1_o_instr_long_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6925_ _0498_ clknet_leaf_50_core_clock dmmu1.page_table\[3\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6856_ _0429_ clknet_leaf_98_core_clock dmmu0.page_table\[1\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5807_ _2808_ _0408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_1968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3999_ _1434_ _1660_ _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6787_ _0360_ clknet_leaf_41_core_clock dmmu1.page_table\[13\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5738_ _2061_ _2760_ _2762_ dmmu1.page_table\[11\]\[3\] _2766_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input81_I c0_sr_bus_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5669_ _2725_ _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_66_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3168__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_10_core_clock clknet_3_1_0_core_clock clknet_leaf_10_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3493__A1 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4690__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output502_I net502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5234__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6959__CLK clknet_leaf_62_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3096__I1 net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4164__I _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4745__A1 _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6339__CLK clknet_leaf_75_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6489__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5473__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3484__A1 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_99_core_clock clknet_3_1_0_core_clock clknet_leaf_99_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3236__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4971_ _2316_ _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3087__I1 net21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4433__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6710_ _0283_ clknet_leaf_26_core_clock dmmu0.page_table\[13\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4984__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3922_ _1368_ _1585_ _1586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3331__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4984__B2 dmmu0.page_table\[14\]\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6641_ _0214_ clknet_leaf_27_core_clock dmmu0.page_table\[15\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3853_ immu_1.page_table\[0\]\[4\] immu_1.page_table\[1\]\[4\] immu_1.page_table\[2\]\[4\]
+ immu_1.page_table\[3\]\[4\] _1409_ _1442_ _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_11_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4736__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5933__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3784_ _1422_ _1427_ _1432_ _1452_ _1453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6572_ _0145_ clknet_leaf_3_core_clock immu_0.page_table\[4\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5523_ _2531_ _2629_ _2631_ dmmu0.page_table\[13\]\[10\] _2643_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_1654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_2030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5454_ _2604_ _0259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput500 net500 c1_i_req_data[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput511 net511 c1_i_req_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput522 net522 dcache_mem_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4405_ _1864_ _1957_ _1959_ net985 _1967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput533 net533 dcache_mem_addr[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5161__A1 _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput544 net544 dcache_mem_i_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5385_ _2563_ _0231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput555 net555 dcache_mem_i_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput566 net566 dcache_wb_i_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput577 net577 dcache_wb_i_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3172__B1 _0921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3711__A2 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7124_ net69 net592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4336_ _1926_ _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput588 net588 ic0_mem_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput599 net599 ic0_mem_ppl_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7055_ net292 net443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4267_ _1861_ _1876_ _1878_ net761 _1885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input233_I dcache_wb_adr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6006_ _2921_ _0494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3218_ _0964_ _0965_ _0842_ _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4198_ _1831_ _1832_ _1833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4672__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3149_ _0898_ _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input400_I inner_wb_i_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3227__A1 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Left_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6908_ _0481_ clknet_leaf_64_core_clock dmmu1.page_table\[5\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3322__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6839_ _0412_ clknet_leaf_44_core_clock dmmu1.page_table\[9\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_1765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3529__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output452_I net452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_2038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6631__CLK clknet_leaf_35_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold280 immu_0.page_table\[8\]\[10\] net1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold291 immu_1.page_table\[5\]\[10\] net1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4159__I net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_2294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6781__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4966__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4718__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4194__A2 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5654__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5694__A2 _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5170_ _2267_ _2430_ _2432_ net774 _2435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4121_ _1306_ _1302_ _0816_ net641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_23_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5446__A2 net379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4052_ _1708_ _1711_ _1712_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3457__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 c0_o_icache_flush net4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4954_ _2273_ _2299_ _2302_ dmmu0.page_table\[7\]\[5\] _2308_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6504__CLK clknet_leaf_8_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3905_ _1385_ immu_0.page_table\[8\]\[5\] _1570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6159__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4885_ _1779_ _1972_ _2259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_7_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6624_ _0197_ clknet_leaf_9_core_clock immu_0.page_table\[0\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3836_ _1408_ _1501_ _1502_ _1503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_12_1973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5382__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3767_ immu_1.page_table\[0\]\[1\] immu_1.page_table\[1\]\[1\] immu_1.page_table\[8\]\[1\]
+ immu_1.page_table\[9\]\[1\] _1435_ _1415_ _1436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6555_ _0128_ clknet_leaf_18_core_clock immu_0.page_table\[6\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3148__I _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6654__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input183_I c1_sr_bus_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5506_ _2634_ _0281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6486_ _0059_ clknet_leaf_33_core_clock dmmu0.page_table\[7\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3698_ _1367_ _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_14_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5437_ _2593_ _0253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input350_I ic1_mem_data[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5368_ _2300_ _2552_ _2554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input44_I c0_o_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4893__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7107_ net398 net575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4319_ _1852_ _1911_ _1914_ immu_1.page_table\[2\]\[3\] _1918_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5299_ net104 _2502_ _2504_ immu_0.page_table\[0\]\[9\] _2513_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_74_2101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7038_ net305 net456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_1108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3448__A1 net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_2_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4948__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_2481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_2492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_2356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_0_core_clock clknet_3_0_0_core_clock clknet_leaf_0_core_clock vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4479__A3 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5676__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3687__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_107_core_clock clknet_3_0_0_core_clock clknet_leaf_107_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_44_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5428__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3439__A1 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__A3 _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6527__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_2095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5061__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3298__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5600__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3611__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6677__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4670_ _2065_ _2123_ _2125_ net1001 _2131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_56_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3621_ _1308_ net267 _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_42_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5364__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3552_ net138 net33 _1267_ _1276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6340_ _0722_ clknet_leaf_74_core_clock immu_1.page_table\[14\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6271_ _0653_ clknet_leaf_89_core_clock immu_1.page_table\[6\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5116__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3483_ _0875_ _1221_ _1222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_45_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5222_ _2467_ _0164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5153_ _2277_ _2414_ _2416_ net894 _2424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_36_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4104_ _1758_ _1759_ _1760_ net701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5084_ _2383_ _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_58_1439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4035_ net107 _1685_ _1695_ _1696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_49_1668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5986_ _2911_ _0484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4937_ _1778_ net84 _2296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_34_1494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input398_I inner_wb_i_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_20 net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4868_ _1809_ _2242_ _2244_ dmmu0.page_table\[9\]\[5\] _2250_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6607_ _0180_ clknet_leaf_5_core_clock immu_0.page_table\[1\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3819_ immu_0.page_table\[0\]\[3\] immu_0.page_table\[1\]\[3\] immu_0.page_table\[2\]\[3\]
+ immu_0.page_table\[3\]\[3\] _1424_ _1455_ _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_69_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4799_ _2209_ _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_15_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6538_ _0111_ clknet_leaf_7_core_clock immu_0.page_table\[7\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6469_ _0042_ clknet_leaf_14_core_clock dmmu0.page_table\[8\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3669__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3542__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6083__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3516__S1 net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5291__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5830__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3841__A1 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5043__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_40_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_2035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_2046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5594__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4397__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4172__I _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5346__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4149__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_2554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5897__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_2418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_2429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4321__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4609__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4085__A1 net11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5282__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5840_ _1808_ _2819_ _2821_ dmmu0.page_table\[1\]\[5\] _2827_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_1281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ _1851_ _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_44_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3200__B _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _1803_ _2157_ _2159_ immu_0.page_table\[15\]\[3\] _2163_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_20_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4653_ _2120_ _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput40 c0_o_mem_data[5] net40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3604_ inner_wb_arbiter.o_sel_sig _1304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
Xinput51 c0_o_mem_high_addr[6] net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3899__A1 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput62 c0_o_req_addr[12] net62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_0_1790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4584_ _2080_ _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_57_1904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput73 c0_o_req_addr[8] net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_57_1915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput84 c0_sr_bus_addr[2] net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_3_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_2019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput95 c0_sr_bus_data_o[12] net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6323_ _0705_ clknet_leaf_70_core_clock dmmu1.page_table\[14\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_1926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3535_ _0840_ _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_29_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3994__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6254_ _0636_ clknet_leaf_84_core_clock immu_1.page_table\[5\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3466_ dmmu1.page_table\[12\]\[11\] dmmu1.page_table\[13\]\[11\] dmmu1.page_table\[14\]\[11\]
+ dmmu1.page_table\[15\]\[11\] _0898_ _0901_ _1205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_0_883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5205_ _1805_ _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_1162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6185_ dmmu1.long_off_reg\[7\] _1864_ _3016_ _3024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3397_ net106 net158 _0884_ _1138_ _1139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_4_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input146_I c1_o_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5136_ _2413_ _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_4_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6065__A2 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5067_ _2271_ _2367_ _2369_ net1036 _2374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5273__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6842__CLK clknet_leaf_67_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input313_I ic0_wb_adr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5812__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4018_ _1654_ _1664_ _1669_ _1679_ _1680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3823__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5025__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4379__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6992__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5969_ _2847_ _2890_ _2892_ net941 _2901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3051__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__CLK clknet_leaf_83_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4000__A1 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3434__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6372__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4839__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output532_I net532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4303__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3106__A3 net52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput400 inner_wb_i_dat[5] net400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_25_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_2211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_67_2222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4067__A1 net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_2233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3814__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_2065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3042__A2 net559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5319__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6715__CLK clknet_leaf_23_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold109 dmmu1.page_table\[11\]\[10\] net843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_65_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4542__A2 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5662__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3320_ dmmu1.page_table\[4\]\[6\] dmmu1.page_table\[5\]\[6\] dmmu1.page_table\[6\]\[6\]
+ dmmu1.page_table\[7\]\[6\] _0888_ _0910_ _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_0_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3750__B1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3251_ _0908_ dmmu1.page_table\[0\]\[4\] _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_33_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6865__CLK clknet_leaf_42_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3182_ _0901_ _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6047__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4058__A1 _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5255__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6941_ _0514_ clknet_leaf_56_core_clock dmmu1.page_table\[2\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3805__A1 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6872_ _0445_ clknet_leaf_52_core_clock dmmu1.page_table\[7\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5007__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5823_ _2816_ _0416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6245__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5754_ _2047_ _2759_ _2761_ net862 _2774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3865__B _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4705_ _2151_ _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5685_ _2735_ _0359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4636_ _2057_ _2108_ _2110_ net861 _2112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6395__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_2094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4533__A2 _2032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5730__A1 _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4567_ _2069_ _2053_ _2055_ net865 _2070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_31_Left_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input263_I dcache_wb_o_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6306_ _0688_ clknet_leaf_89_core_clock immu_1.page_table\[3\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3518_ dmmu1.page_table\[12\]\[12\] dmmu1.page_table\[13\]\[12\] dmmu1.page_table\[14\]\[12\]
+ dmmu1.page_table\[15\]\[12\] _0886_ net121 _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4498_ _2024_ _0692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6237_ _0619_ clknet_leaf_87_core_clock immu_1.page_table\[2\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3449_ net154 dmmu1.long_off_reg\[4\] _1189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4297__A1 _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6168_ _1764_ _1767_ _3014_ _0563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5119_ _2404_ _0124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4049__A1 net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5246__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6099_ _1891_ _1892_ _2030_ _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_20_1891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_40_Left_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5549__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4221__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4221__B2 immu_1.page_table\[9\]\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6738__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4772__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4450__I net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3407__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3958__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6888__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5485__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput230 dcache_wb_4_burst net230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput241 dcache_wb_adr[19] net241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput252 dcache_wb_adr[7] net252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6029__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput263 dcache_wb_o_dat[1] net263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput274 dcache_wb_stb net274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput285 ic0_mem_data[17] net285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput296 ic0_mem_data[27] net296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_89_core_clock clknet_3_4_0_core_clock clknet_leaf_89_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5788__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3894__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4763__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5470_ _2612_ _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4421_ _1978_ _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput704 net704 inner_wb_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4515__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5712__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7140_ net389 net604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4352_ _1936_ _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3303_ _0897_ _1047_ _0912_ _1048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7071_ net353 net506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4283_ _1895_ _1893_ _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3234_ dmmu1.page_table\[0\]\[3\] dmmu1.page_table\[1\]\[3\] dmmu1.page_table\[2\]\[3\]
+ dmmu1.page_table\[3\]\[3\] _0899_ _0902_ _0981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6022_ _2931_ _0500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3165_ net123 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5228__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3096_ net130 net25 _0850_ _0851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4535__I net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6924_ _0497_ clknet_leaf_53_core_clock dmmu1.page_table\[3\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4451__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input109_I c1_o_icache_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6855_ _0428_ clknet_leaf_97_core_clock dmmu0.page_table\[1\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5806_ _2786_ _2802_ _2804_ dmmu1.page_table\[9\]\[3\] _2808_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4203__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6786_ _0359_ clknet_leaf_43_core_clock dmmu1.page_table\[13\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3998_ immu_1.page_table\[12\]\[8\] immu_1.page_table\[13\]\[8\] immu_1.page_table\[14\]\[8\]
+ immu_1.page_table\[15\]\[8\] _1441_ _1540_ _1660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_17_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5737_ _2765_ _0381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5951__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3087__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input380_I ic1_wb_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5668_ _1828_ _2028_ _2031_ _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_5_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input74_I c0_o_req_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4619_ _2069_ _2090_ _2092_ immu_1.page_table\[13\]\[7\] _2100_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5599_ _2687_ _0321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6410__CLK clknet_leaf_109_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3550__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5219__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4690__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3493__A2 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_1740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3876__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3556__I0 net140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5170__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3181__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6903__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4970_ _1977_ _2173_ _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__3236__A2 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4433__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5630__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3921_ immu_0.page_table\[0\]\[6\] immu_0.page_table\[1\]\[6\] immu_0.page_table\[2\]\[6\]
+ immu_0.page_table\[3\]\[6\] _1424_ _1455_ _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_50_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4984__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6640_ _0213_ clknet_leaf_25_core_clock dmmu0.page_table\[15\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3852_ immu_1.page_table\[8\]\[4\] immu_1.page_table\[9\]\[4\] immu_1.page_table\[10\]\[4\]
+ immu_1.page_table\[11\]\[4\] _1409_ _1442_ _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_6_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5933__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__A2 _2156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6571_ _0144_ clknet_leaf_6_core_clock immu_0.page_table\[4\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3783_ _1433_ _1438_ _1451_ _0813_ _1452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_41_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5522_ _2642_ _0289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5453_ immu_1.high_addr_off\[0\] _1824_ _2603_ _2604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput501 net501 c1_i_req_data[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4044__S0 _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput512 net512 c1_i_req_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput523 net523 dcache_mem_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4404_ _1966_ _0656_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput534 net534 dcache_mem_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_1953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput545 net545 dcache_mem_i_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_22_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5384_ _2463_ _2553_ _2555_ dmmu0.page_table\[11\]\[7\] _2563_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput556 net556 dcache_mem_i_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3172__A1 _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput567 net567 dcache_wb_i_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3172__B2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7123_ net68 net591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput578 net578 dcache_wb_i_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4335_ _1828_ _1839_ _1873_ _1926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xoutput589 net589 ic0_mem_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3711__A3 net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6433__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7054_ net291 net442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4266_ _1884_ _0600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6005_ net199 _2906_ _2908_ dmmu1.page_table\[4\]\[11\] _2921_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3217_ _0897_ _0895_ _0965_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3370__S _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4197_ net185 net184 net183 net182 _1832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__4672__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input226_I dcache_mem_o_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6583__CLK clknet_leaf_21_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3148_ _0886_ _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_55_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3079_ _0840_ _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__3227__A2 _0973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3858__S0 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6907_ _0480_ clknet_leaf_63_core_clock dmmu1.page_table\[5\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _0411_ clknet_leaf_49_core_clock dmmu1.page_table\[9\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4027__I1 _1687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_45_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6769_ _0342_ clknet_leaf_39_core_clock dmmu0.page_table\[5\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3538__I0 net146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5688__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3163__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold270 immu_1.page_table\[7\]\[5\] net1004 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_output445_I net445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold281 immu_1.page_table\[8\]\[2\] net1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold292 immu_1.page_table\[4\]\[4\] net1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6101__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_2295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5860__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4415__A1 _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_1289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3849__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5612__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4966__A2 _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6306__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4718__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5915__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_2097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3963__B _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4026__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3455__S _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6456__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3529__I0 net142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5143__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3154__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4120_ _1306_ _1302_ _0815_ net640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_78_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4051_ _1699_ _1709_ _1710_ _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_53_1792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3190__S _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4654__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 c0_o_instr_long_addr[0] net5 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_2008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4953_ _2307_ _0055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3904_ _1391_ _1567_ _1568_ _1569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_30_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3857__C _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6159__A1 _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4884_ _1776_ _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_69_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6623_ _0196_ clknet_leaf_6_core_clock immu_0.page_table\[0\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3835_ _1415_ _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_7_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6554_ _0127_ clknet_leaf_19_core_clock immu_0.page_table\[6\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3766_ _1409_ _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5382__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5505_ _2451_ _2630_ _2632_ dmmu0.page_table\[13\]\[1\] _2634_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3393__A1 _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6485_ _0058_ clknet_leaf_26_core_clock dmmu0.page_table\[7\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3697_ _1366_ _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_14_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input176_I c1_o_req_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5436_ _2527_ _2582_ _2584_ net834 _2593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6949__CLK clknet_leaf_53_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3145__A1 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5367_ _2552_ _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_input343_I ic1_mem_data[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4893__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7106_ net397 net574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4318_ _1917_ _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5298_ _2512_ _0195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input37_I c0_o_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7037_ net304 net455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4249_ _1872_ net189 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__5842__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6329__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4948__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_1_0_core_clock clknet_0_core_clock clknet_3_1_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_4_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3783__B _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3384__A1 net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4581__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4008__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_2493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6173__I1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_2368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3687__A2 net364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4636__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_2006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5061__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3298__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3611__A2 net256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_78_Left_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3620_ _1313_ net695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_42_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5364__A2 _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3693__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3551_ _1275_ net546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6270_ _0652_ clknet_leaf_88_core_clock immu_1.page_table\[6\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5116__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_2012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3482_ dmmu0.page_table\[12\]\[11\] dmmu0.page_table\[13\]\[11\] dmmu0.page_table\[14\]\[11\]
+ dmmu0.page_table\[15\]\[11\] _0863_ _0866_ _1221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_62_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5221_ _2332_ _2446_ _2448_ net892 _2467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_59_1990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5152_ _2423_ _0138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6077__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4103_ _1535_ net272 _1760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3712__I _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5083_ _2140_ _2381_ _2383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4034_ _0813_ _1694_ _1695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5985_ _2782_ _2907_ _2909_ dmmu1.page_table\[4\]\[1\] _2911_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_2016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6621__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4936_ _2294_ _2295_ _1771_ _0050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_10 net392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_21 net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3159__I _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4867_ _2249_ _0027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6001__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input293_I ic0_mem_data[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6606_ _0179_ clknet_leaf_15_core_clock immu_0.page_table\[1\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3818_ _1485_ net665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4798_ _2140_ _2207_ _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3366__A1 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6771__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6537_ _0110_ clknet_leaf_4_core_clock immu_0.page_table\[7\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3749_ _1405_ _1408_ _1418_ _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_28_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6468_ _0041_ clknet_leaf_22_core_clock dmmu0.page_table\[8\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4315__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5419_ _2583_ _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6399_ _0781_ clknet_leaf_108_core_clock immu_0.page_table\[15\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3669__A2 net375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5291__A1 _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_2172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5043__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_2047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5594__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5346__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3357__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_2419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3747__I3 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3109__A1 net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6059__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3532__I _1265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4609__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5806__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6644__CLK clknet_leaf_35_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5770_ _2785_ _0394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_44_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A2 _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6794__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4721_ _2162_ _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4652_ _2103_ _2108_ _2110_ immu_1.page_table\[12\]\[9\] _2120_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3348__A1 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3603_ _1302_ net382 _1303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput30 c0_o_mem_data[10] net30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput41 c0_o_mem_data[6] net41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput52 c0_o_mem_high_addr[7] net52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4583_ _2059_ _2075_ _2077_ immu_1.page_table\[14\]\[2\] _2080_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput63 c0_o_req_addr[13] net63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_80_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput74 c0_o_req_addr[9] net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6322_ _0704_ clknet_leaf_70_core_clock dmmu1.page_table\[14\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3534_ _1266_ net553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput85 c0_sr_bus_addr[3] net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_57_1927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput96 c0_sr_bus_data_o[1] net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6253_ _0635_ clknet_leaf_83_core_clock immu_1.page_table\[5\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3465_ _0841_ _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_38_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5204_ _2456_ _0157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6184_ _3023_ _0570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3396_ _0894_ _1128_ _1137_ _1138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3520__A1 net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5135_ _1789_ _2412_ _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4538__I net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input139_I c1_o_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5066_ _2373_ _0102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5273__A1 net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4017_ _1301_ _1678_ _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3823__A2 _1489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input306_I ic0_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5025__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5369__I _2554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5968_ _2900_ _0477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3587__A1 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4784__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4919_ _1994_ _2260_ _2262_ net778 _2282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5899_ _2786_ _2856_ _2858_ net921 _2862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3434__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6517__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4839__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3106__A4 net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput401 inner_wb_i_dat[6] net401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_60_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output525_I net525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6667__CLK clknet_leaf_103_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_79_core_clock clknet_3_5_0_core_clock clknet_leaf_79_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_67_2212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3814__A2 net705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_2109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_2011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5567__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5319__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4527__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6197__CLK clknet_leaf_1_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A3 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3750__A1 _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3750__B2 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3463__S _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3250_ dmmu1.page_table\[1\]\[4\] _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_24_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3181_ _0915_ _0924_ _0929_ _0895_ _0930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__5255__A1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6940_ _0513_ clknet_leaf_57_core_clock dmmu1.page_table\[2\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6871_ _0444_ clknet_leaf_48_core_clock dmmu1.page_table\[7\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5007__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5822_ _2047_ _2801_ _2803_ dmmu1.page_table\[9\]\[11\] _2816_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_27_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3569__A1 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5753_ _2773_ _0389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4704_ _2101_ _2139_ _2142_ immu_1.page_table\[10\]\[8\] _2151_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5684_ _2067_ _2726_ _2728_ net772 _2735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_1517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4635_ _2111_ _0742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4566_ _1863_ _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_69_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6305_ _0687_ clknet_leaf_93_core_clock immu_1.page_table\[3\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3517_ _0905_ _1254_ _1255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4497_ _1864_ _2014_ _2016_ immu_1.page_table\[3\]\[7\] _2024_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input256_I dcache_wb_o_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6236_ _0618_ clknet_leaf_80_core_clock immu_1.page_table\[2\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3448_ net154 dmmu1.long_off_reg\[4\] _1188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4297__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6167_ _1535_ net255 _1895_ _3014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3379_ net47 dmmu0.long_off_reg\[2\] _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5118_ _2269_ _2398_ _2400_ immu_0.page_table\[6\]\[3\] _2404_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6098_ _2973_ _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_38_1619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5246__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5049_ _2328_ _2352_ _2354_ immu_0.page_table\[9\]\[8\] _2363_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3352__S0 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5549__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_102_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4757__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5827__I _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3548__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4221__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3980__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3407__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5182__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3791__B _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3732__A1 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_52_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput220 dcache_mem_o_data[15] net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3082__I _0843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput231 dcache_wb_adr[0] net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput242 dcache_wb_adr[1] net242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput253 dcache_wb_adr[8] net253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput264 dcache_wb_o_dat[2] net264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput275 dcache_wb_we net275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput286 ic0_mem_data[18] net286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput297 ic0_mem_data[28] net297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5788__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_1517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3799__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3894__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6832__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4420_ _1973_ _1977_ _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_1_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5712__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3723__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4351_ _1861_ _1927_ _1929_ net775 _1936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3302_ dmmu1.page_table\[8\]\[5\] dmmu1.page_table\[9\]\[5\] dmmu1.page_table\[10\]\[5\]
+ dmmu1.page_table\[11\]\[5\] _0908_ _0910_ _1047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_7070_ net342 net495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4282_ _1769_ _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XANTENNA__6982__CLK clknet_leaf_73_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6021_ _2788_ _2924_ _2926_ dmmu1.page_table\[3\]\[4\] _2931_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3233_ dmmu1.page_table\[4\]\[3\] dmmu1.page_table\[5\]\[3\] dmmu1.page_table\[6\]\[3\]
+ dmmu1.page_table\[7\]\[3\] _0899_ _0902_ _0980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_20_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3164_ _0904_ _0913_ _0895_ _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_20_1166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5228__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6212__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3095_ _0840_ _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_59_1387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _0496_ clknet_leaf_53_core_clock dmmu1.page_table\[3\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4451__A2 _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _0427_ clknet_leaf_37_core_clock dmmu0.page_table\[1\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6362__CLK clknet_leaf_75_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5805_ _2807_ _0407_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6785_ _0358_ clknet_leaf_49_core_clock dmmu1.page_table\[13\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4203__A2 _1834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3997_ _1440_ _1658_ _1659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4551__I _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5736_ _2059_ _2760_ _2762_ dmmu1.page_table\[11\]\[2\] _2765_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5951__A2 _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_6_0_core_clock clknet_0_core_clock clknet_3_6_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_66_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3962__A1 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5667_ _2724_ _0352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input373_I ic1_wb_adr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4618_ _2099_ _0737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5598_ _2453_ _2681_ _2684_ net903 _2687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4506__A3 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input67_I c0_o_req_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4911__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4549_ _2057_ _2053_ _2055_ net812 _2058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6219_ _0601_ clknet_leaf_87_core_clock immu_1.page_table\[7\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_2019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5219__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4690__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7102__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4978__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6705__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3876__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output592_I net592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5155__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3556__I1 net35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6235__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6385__CLK clknet_leaf_72_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4433__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3920_ _1375_ _1583_ _1584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3851_ _1515_ _1516_ _1446_ _1517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5394__B1 _2554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6570_ _0143_ clknet_leaf_17_core_clock immu_0.page_table\[4\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3782_ net705 _1447_ _1450_ _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5933__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3944__A1 net112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5521_ _2529_ _2630_ _2632_ net1092 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5452_ _2602_ _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_2_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput502 net502 c1_i_req_data[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4044__S1 _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_2092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4403_ _1861_ _1957_ _1959_ net937 _1966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput513 net513 c1_i_req_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput524 net524 dcache_mem_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5383_ _2562_ _0230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_65_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput535 net535 dcache_mem_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput546 net546 dcache_mem_i_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput557 net557 dcache_mem_i_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7122_ net67 net590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput568 net568 dcache_wb_i_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4334_ _1925_ _0627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput579 net579 dcache_wb_i_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_5_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5449__A1 net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7053_ net290 net441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4265_ _1858_ _1876_ _1878_ net1004 _1884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4121__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6004_ _2920_ _0493_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3216_ _0962_ _0963_ _0912_ _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4196_ net187 net186 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4672__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3147_ _0896_ _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_input121_I c1_o_mem_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input219_I dcache_mem_o_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3078_ _0819_ _0820_ _0840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_49_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3858__S1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6906_ _0479_ clknet_leaf_60_core_clock dmmu1.page_table\[5\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6878__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6837_ _0410_ clknet_leaf_48_core_clock dmmu1.page_table\[9\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3098__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6768_ _0341_ clknet_leaf_40_core_clock dmmu0.page_table\[5\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3935__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5719_ _2754_ _0374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_66_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6699_ _0272_ clknet_leaf_30_core_clock dmmu0.page_table\[4\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_1491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5688__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3538__I1 net41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6258__CLK clknet_leaf_84_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold260 dmmu0.page_table\[14\]\[1\] net994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3163__A2 _0911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold271 immu_1.page_table\[11\]\[9\] net1005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold282 immu_0.page_table\[13\]\[0\] net1016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold293 immu_0.page_table\[15\]\[10\] net1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_output438_I net438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6101__A2 _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_2296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5860__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4415__A2 _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5612__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__I1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3849__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5376__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5128__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3963__C _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4026__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3529__I1 net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4351__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4103__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4050_ net10 immu_0.high_addr_off\[5\] _1710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_21_1250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_1793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput6 c0_o_instr_long_addr[1] net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4952_ _2271_ _2299_ _2302_ dmmu0.page_table\[7\]\[4\] _2307_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3903_ _1463_ immu_0.page_table\[11\]\[5\] _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4883_ _2257_ _0035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6159__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3834_ _1499_ _1500_ _1439_ _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6622_ _0195_ clknet_leaf_16_core_clock immu_0.page_table\[0\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6553_ _0126_ clknet_leaf_19_core_clock immu_0.page_table\[6\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3765_ _1416_ _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_12_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6400__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5504_ _2633_ _0280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6484_ _0057_ clknet_leaf_13_core_clock dmmu0.page_table\[7\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3696_ net314 _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_28_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5435_ _2592_ _0252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3145__A2 net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input169_I c1_o_req_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ _1781_ _1977_ _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_61_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6550__CLK clknet_leaf_3_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4893__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7105_ net396 net573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4317_ _1849_ _1911_ _1914_ net848 _1917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5297_ net103 _2502_ _2504_ immu_0.page_table\[0\]\[8\] _2512_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6095__A1 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7036_ net303 net454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input336_I ic1_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4248_ net190 _1872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__5842__A1 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4179_ net103 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5358__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_14_Right_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3556__S _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3783__C _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4581__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4008__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_2494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4333__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3767__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_2369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_23_Right_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4636__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3090__I _0847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_2075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5061__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3072__A1 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Right_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6423__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3550_ net137 net32 _1267_ _1275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_1984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6573__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3481_ dmmu0.page_table\[8\]\[11\] dmmu0.page_table\[9\]\[11\] dmmu0.page_table\[10\]\[11\]
+ dmmu0.page_table\[11\]\[11\] _0871_ _0867_ _1220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_11_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5220_ _2466_ _0163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_59_1980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_41_Right_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5521__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5151_ _2275_ _2414_ _2416_ immu_0.page_table\[5\]\[6\] _2423_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6077__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4102_ _1350_ net326 _1360_ _1759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5082_ _2381_ _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_36_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5824__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ _1502_ _1688_ _1693_ net705 _1694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_75_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__I _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3868__C _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_50_Right_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5984_ _2910_ _0483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4935_ _1796_ _2290_ _2291_ _1845_ _2295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_11 net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_22 net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4866_ _1806_ _2242_ _2244_ dmmu0.page_table\[9\]\[4\] _2249_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6001__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6916__CLK clknet_leaf_54_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_107_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6605_ _0178_ clknet_leaf_15_core_clock immu_0.page_table\[1\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_1559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3817_ net236 _1484_ _1360_ _1485_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4797_ _2207_ _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_55_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input286_I ic0_mem_data[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3748_ _1408_ _1417_ _1418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6536_ _0109_ clknet_leaf_100_core_clock immu_0.page_table\[8\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3679_ _1348_ net377 _1353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6467_ _0040_ clknet_leaf_28_core_clock dmmu0.page_table\[8\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4315__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5418_ _2300_ _2581_ _2583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6398_ _0780_ clknet_leaf_108_core_clock immu_0.page_table\[15\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4866__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5349_ _2543_ _0215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_69_core_clock clknet_3_4_0_core_clock clknet_leaf_69_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5666__I1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_57_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5291__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3921__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6446__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3778__C _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5579__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7110__I net401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_2162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5043__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_2173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_2051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_2037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_2048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6596__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5503__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5806__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4609__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5282__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3293__A1 _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3045__A1 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ _1800_ _2157_ _2159_ immu_0.page_table\[15\]\[2\] _2162_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_29_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ _2119_ _0750_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput20 c0_o_mem_addr[1] net20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3602_ _1301_ _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput31 c0_o_mem_data[11] net31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5742__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3979__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4582_ _2079_ _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput42 c0_o_mem_data[7] net42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput53 c0_o_mem_long_mode net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_12_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput64 c0_o_req_addr[14] net64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput75 c0_o_req_ppl_submit net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3533_ net144 net39 _0850_ _1266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6321_ _0703_ clknet_leaf_96_core_clock dmmu1.page_table\[14\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_1906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput86 c0_sr_bus_addr[4] net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput97 c0_sr_bus_data_o[2] net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6252_ _0634_ clknet_leaf_88_core_clock immu_1.page_table\[5\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3464_ _1203_ net531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6319__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5203_ _2455_ _2447_ _2449_ net939 _2456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6183_ dmmu1.long_off_reg\[6\] _1861_ _3016_ _3023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3395_ _0915_ _1131_ _1136_ _0894_ _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_58_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5134_ _2205_ _2296_ _2412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6469__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5065_ _2269_ _2367_ _2369_ net971 _2373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4016_ _1378_ _1672_ _1677_ _1381_ _1678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__5273__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3284__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4554__I _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input201_I c1_sr_bus_data_o[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5025__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3036__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5967_ _2794_ _2890_ _2892_ net1077 _2900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3587__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4784__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4918_ _2281_ _0046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5898_ _2861_ _0446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_2068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input97_I c0_sr_bus_data_o[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4849_ _1994_ _2223_ _2225_ net965 _2238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4536__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6519_ _0092_ clknet_leaf_109_core_clock immu_0.page_table\[9\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_1654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3834__S _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4839__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7105__I net396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput402 inner_wb_i_dat[7] net402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_76_1338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_2213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3275__A1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_1073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_14_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4527__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4527__B2 dmmu1.page_table\[14\]\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3750__A2 _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3543__I _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6611__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3180_ _0926_ _0928_ _0915_ _0929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_20_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5255__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6761__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3266__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4463__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _0443_ clknet_leaf_67_core_clock dmmu1.page_table\[8\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5007__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5821_ _2815_ _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_27_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3569__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5963__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5752_ _2105_ _2759_ _2761_ net843 _2773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_56_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4703_ _2150_ _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5683_ _2734_ _0358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4634_ _2051_ _2108_ _2110_ net907 _2111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4565_ _2068_ _0715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3881__C _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6304_ _0686_ clknet_leaf_80_core_clock immu_1.page_table\[3\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3516_ dmmu1.page_table\[8\]\[12\] dmmu1.page_table\[9\]\[12\] dmmu1.page_table\[10\]\[12\]
+ dmmu1.page_table\[11\]\[12\] _0886_ net121 _1254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4496_ _2023_ _0691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_4_Right_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6235_ _0617_ clknet_leaf_81_core_clock immu_1.page_table\[2\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6291__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3447_ net155 dmmu1.long_off_reg\[5\] _1187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input151_I c1_o_mem_high_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input249_I dcache_wb_adr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3344__I2 dmmu1.page_table\[14\]\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3378_ net47 dmmu0.long_off_reg\[2\] _1120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6166_ _3013_ _0562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5117_ _2403_ _0123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6097_ net200 _2957_ _2959_ dmmu1.page_table\[1\]\[12\] _2973_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5246__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5048_ _2362_ _0095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3257__A1 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input12_I c0_o_instr_long_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3352__S1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6999_ _0572_ clknet_leaf_103_core_clock icore_sregs.c1_disable vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_24_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4757__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_2076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4509__A1 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5706__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5182__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6634__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3732__A2 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output635_I net635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5485__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput210 c1_sr_bus_we net210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3496__A1 net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6784__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput221 dcache_mem_o_data[1] net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput232 dcache_wb_adr[10] net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput243 dcache_wb_adr[20] net243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput254 dcache_wb_adr[9] net254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput265 dcache_wb_o_dat[3] net265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput276 ic0_mem_ack net276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput287 ic0_mem_data[19] net287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput298 ic0_mem_data[29] net298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3248__A1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3799__A2 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4350_ _1935_ _0633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3301_ _0907_ _1045_ _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4281_ _1893_ _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_39_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6020_ _2930_ _0499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3232_ _0977_ _0978_ _0884_ _0979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_20_1101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3487__A1 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I c0_o_icache_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3163_ _0907_ _0911_ _0912_ _0913_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5228__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3094_ _0849_ net537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3222__B _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6922_ _0495_ clknet_leaf_63_core_clock dmmu1.page_table\[4\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6507__CLK clknet_leaf_8_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6853_ _0426_ clknet_leaf_41_core_clock dmmu0.page_table\[1\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5804_ _2784_ _2802_ _2804_ dmmu1.page_table\[9\]\[2\] _2807_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6784_ _0357_ clknet_leaf_44_core_clock dmmu1.page_table\[13\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3996_ immu_1.page_table\[8\]\[8\] immu_1.page_table\[9\]\[8\] immu_1.page_table\[10\]\[8\]
+ immu_1.page_table\[11\]\[8\] _1441_ _1540_ _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_29_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5735_ _2764_ _0380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_50_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6657__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input199_I c1_sr_bus_data_o[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5666_ dmmu0.long_off_reg\[7\] _1815_ _2716_ _2724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5164__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4617_ _2067_ _2090_ _2092_ net1064 _2099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5597_ _2686_ _0320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input366_I ic1_wb_adr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4911__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4548_ _1845_ _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_44_1635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6113__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3183__I net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4479_ _1838_ _1874_ _1891_ _2013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_22_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6218_ _0600_ clknet_leaf_85_core_clock immu_1.page_table\[7\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3478__A1 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6149_ _1848_ _3000_ _3002_ net1015 _3005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5219__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4427__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4978__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3650__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4742__I _2174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5927__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output585_I net585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3402__A1 net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5155__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4189__I _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3308__I2 dmmu0.page_table\[14\]\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3469__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4666__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3641__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3850_ immu_1.page_table\[4\]\[4\] immu_1.page_table\[5\]\[4\] immu_1.page_table\[6\]\[4\]
+ immu_1.page_table\[7\]\[4\] _1441_ _1442_ _1516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3781_ _1440_ _1448_ _1449_ _1444_ _1415_ _1450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__5394__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3268__I net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _2641_ _0288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5451_ _1834_ _2601_ _2602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_2082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4402_ _1965_ _0655_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput503 net503 c1_i_req_data[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput514 net514 c1_i_req_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_2055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput525 net525 dcache_mem_addr[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5382_ _2461_ _2553_ _2555_ dmmu0.page_table\[11\]\[6\] _2562_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput536 net536 dcache_mem_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_61_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput547 net547 dcache_mem_i_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7121_ net66 net589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput558 net558 dcache_mem_i_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4333_ _1870_ _1910_ _1913_ immu_1.page_table\[2\]\[10\] _1925_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput569 net569 dcache_wb_i_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5449__A2 _1836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4264_ _1883_ _0599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7052_ net289 net440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3215_ dmmu1.page_table\[8\]\[2\] dmmu1.page_table\[9\]\[2\] dmmu1.page_table\[10\]\[2\]
+ dmmu1.page_table\[11\]\[2\] _0899_ _0902_ _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6003_ _2851_ _2906_ _2908_ net970 _2920_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4121__A2 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4195_ net195 _1830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_19_Left_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_1715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3146_ net122 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_39_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4409__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3880__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3077_ _0839_ net473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_1038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_2015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input114_I c1_o_instr_long_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6905_ _0478_ clknet_leaf_59_core_clock dmmu1.page_table\[5\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6836_ _0409_ clknet_leaf_48_core_clock dmmu1.page_table\[9\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5909__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6767_ _0340_ clknet_leaf_46_core_clock dmmu0.page_table\[5\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3979_ immu_0.page_table\[8\]\[7\] immu_0.page_table\[9\]\[7\] immu_0.page_table\[10\]\[7\]
+ immu_0.page_table\[11\]\[7\] _1487_ _1390_ _1642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5718_ _2101_ _2743_ _2745_ net1065 _2754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6698_ _0271_ clknet_leaf_31_core_clock dmmu0.page_table\[4\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5137__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5649_ _2714_ _0344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5688__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4896__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold250 dmmu1.page_table\[2\]\[8\] net984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold261 dmmu0.page_table\[14\]\[12\] net995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold272 immu_1.page_table\[7\]\[0\] net1006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold283 dmmu0.page_table\[12\]\[0\] net1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold294 dmmu0.page_table\[6\]\[8\] net1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_2297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7113__I net404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5860__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3871__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output500_I net500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5073__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5612__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3623__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5376__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6972__CLK clknet_leaf_62_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3088__I _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3482__S0 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_64_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5128__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6202__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3234__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6352__CLK clknet_leaf_71_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4103__A2 net272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3551__I _1275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 c0_o_instr_long_addr[2] net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ _2306_ _0054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3902_ _1385_ immu_0.page_table\[10\]\[5\] _1567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_1656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4882_ _1996_ _2241_ _2243_ net883 _2257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6621_ _0194_ clknet_leaf_15_core_clock immu_0.page_table\[0\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3833_ immu_1.page_table\[0\]\[3\] immu_1.page_table\[1\]\[3\] immu_1.page_table\[2\]\[3\]
+ immu_1.page_table\[3\]\[3\] _1435_ _1469_ _1500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_7_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6552_ _0125_ clknet_leaf_4_core_clock immu_0.page_table\[6\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3764_ _1410_ _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3473__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5503_ _2444_ _2630_ _2632_ dmmu0.page_table\[13\]\[0\] _2633_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_6_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6483_ _0056_ clknet_leaf_29_core_clock dmmu0.page_table\[7\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3726__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3695_ _1363_ _1364_ _1365_ net662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_67_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5434_ _2463_ _2582_ _2584_ net814 _2592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_1610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3225__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4878__B1 _2243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5365_ _2551_ _0223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7104_ net389 net566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4316_ _1916_ _0618_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5296_ _2511_ _0194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6095__A2 _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4557__I _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7035_ net302 net453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_59_core_clock clknet_3_7_0_core_clock clknet_leaf_59_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4247_ _1871_ _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6845__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input231_I dcache_wb_adr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input329_I ic0_wb_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5842__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4178_ _1816_ _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_2_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3129_ _0878_ _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_2_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6995__CLK clknet_leaf_95_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4802__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_2090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6819_ _0392_ clknet_leaf_47_core_clock dmmu1.page_table\[10\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5358__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6225__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4581__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7108__I net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_98_core_clock clknet_3_1_0_core_clock clknet_leaf_98_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_76_2484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6375__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_2495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output450_I net450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_2359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3767__S1 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4097__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3844__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3072__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4021__A1 net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6718__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3480_ _0841_ _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_62_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5521__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6868__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5150_ _2422_ _0137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_55_1867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6077__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4101_ _1348_ net380 _1758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5081_ _1790_ _2297_ _2381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_36_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4088__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5285__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4032_ _1415_ _1690_ _1692_ _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_47_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5037__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5983_ _2776_ _2907_ _2909_ dmmu1.page_table\[4\]\[0\] _2910_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6248__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4934_ net407 _2293_ _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4045__C _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4865_ _2248_ _0026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_12 net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_23 _1268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6001__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6604_ _0177_ clknet_leaf_7_core_clock immu_0.page_table\[1\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3816_ _1422_ _1459_ _1468_ _1473_ _1483_ _1484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_74_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4012__A1 _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6398__CLK clknet_leaf_108_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ _1790_ _2206_ _2207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6535_ _0108_ clknet_leaf_1_core_clock immu_0.page_table\[8\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3747_ _1411_ _1412_ _1413_ _1414_ _1415_ _1416_ _1417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA_input181_I c1_sr_bus_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input279_I ic0_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6466_ _0039_ clknet_leaf_28_core_clock dmmu0.page_table\[8\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3678_ _1349_ _1351_ _1352_ net681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4315__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5417_ _2581_ _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6397_ _0779_ clknet_leaf_107_core_clock immu_0.page_table\[15\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5348_ _2457_ _2536_ _2538_ dmmu0.page_table\[15\]\[4\] _2543_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input42_I c0_o_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3191__I _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4079__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5279_ _2501_ _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_39_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3826__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3921__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_2163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_2030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_2027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4251__A1 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_2038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_2049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_2085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output498_I net498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_78_2535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5200__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_2546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output665_I net665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_2557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5503__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5267__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5806__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_2007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5019__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3045__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6540__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4650_ _2101_ _2108_ _2110_ immu_1.page_table\[12\]\[8\] _2119_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_1069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3601_ icache_arbiter.o_sel_sig _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
Xinput10 c0_o_instr_long_addr[5] net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5742__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput21 c0_o_mem_addr[2] net21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 c0_o_mem_data[12] net32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3979__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4581_ _2057_ _2075_ _2077_ immu_1.page_table\[14\]\[1\] _2079_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput43 c0_o_mem_data[8] net43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6690__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput54 c0_o_mem_req net54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6320_ _0702_ clknet_leaf_69_core_clock dmmu1.page_table\[14\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3532_ _1265_ net552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput65 c0_o_req_addr[15] net65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_57_1907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput76 c0_sr_bus_addr[0] net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_40_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput87 c0_sr_bus_addr[5] net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput98 c0_sr_bus_data_o[3] net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_57_1929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6251_ _0633_ clknet_leaf_85_core_clock immu_1.page_table\[5\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3463_ _1186_ _1202_ _0884_ _1203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5202_ _1802_ _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_0_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6182_ _3022_ _0569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3394_ net123 _1133_ _1135_ _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5133_ _2411_ _0131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_4_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ _2372_ _0101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3808__A1 _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4015_ _1377_ _1674_ _1676_ _1677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4481__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5966_ _2899_ _0476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3036__A2 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5430__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_106_core_clock clknet_3_0_0_core_clock clknet_leaf_106_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4917_ _1821_ _2260_ _2262_ net990 _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4784__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5981__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _2784_ _2856_ _2858_ dmmu1.page_table\[7\]\[2\] _2861_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input396_I inner_wb_i_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4848_ _2237_ _0020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3419__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4536__A2 _2032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ _2197_ _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6518_ _0091_ clknet_leaf_8_core_clock immu_0.page_table\[9\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6449_ _0022_ clknet_leaf_99_core_clock dmmu0.page_table\[10\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3135__B _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput403 inner_wb_i_dat[8] net403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6413__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_2214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7121__I net66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3814__A4 _1481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6563__CLK clknet_leaf_18_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3822__I1 _1488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4527__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5724__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4463__A1 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7031__I net406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3266__A2 _0994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5820_ _2105_ _2801_ _2803_ net917 _2815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5751_ _2772_ _0388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5963__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _2069_ _2139_ _2142_ net754 _2150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5682_ _2065_ _2726_ _2728_ dmmu1.page_table\[13\]\[5\] _2734_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4633_ _2109_ _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_68_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4074__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4564_ _2067_ _2053_ _2055_ net944 _2068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_2086 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6303_ _0685_ clknet_leaf_79_core_clock immu_1.page_table\[3\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3515_ _1251_ _1252_ _0896_ _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6436__CLK clknet_leaf_100_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4495_ _1861_ _2014_ _2016_ immu_1.page_table\[3\]\[6\] _2023_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3734__I net366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5479__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6234_ _0616_ clknet_leaf_93_core_clock immu_1.page_table\[0\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3446_ _1179_ _1185_ _1186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_1563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6165_ _2851_ _2999_ _3001_ immu_1.page_table\[8\]\[10\] _3013_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3377_ net53 _0859_ _1119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_77_1604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input144_I c1_o_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5116_ _2267_ _2398_ _2400_ immu_0.page_table\[6\]\[2\] _2403_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6586__CLK clknet_leaf_21_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6096_ _2972_ _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5047_ _2277_ _2352_ _2354_ net785 _2362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input311_I ic0_wb_adr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6998_ _0571_ clknet_leaf_95_core_clock dmmu1.long_off_reg\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_24_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4757__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5949_ _1828_ _1873_ _2030_ _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_36_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4509__A2 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5706__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5182__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_69_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7116__I net392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6131__A1 net559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6929__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output628_I net628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput200 c1_sr_bus_data_o[12] net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput211 core_reset net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
Xinput222 dcache_mem_o_data[2] net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput233 dcache_wb_adr[11] net233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput244 dcache_wb_adr[21] net244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput255 dcache_wb_cyc net255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput266 dcache_wb_o_dat[4] net266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput277 ic0_mem_data[0] net277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput288 ic0_mem_data[1] net288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput299 ic0_mem_data[2] net299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4445__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5642__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4056__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6459__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3982__C _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3803__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3184__A1 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4381__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3300_ dmmu1.page_table\[12\]\[5\] dmmu1.page_table\[13\]\[5\] dmmu1.page_table\[14\]\[5\]
+ dmmu1.page_table\[15\]\[5\] _0888_ _0910_ _1045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_4280_ _1838_ _1891_ _1892_ _1893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_43_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3231_ _0879_ _0883_ _0978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3162_ net123 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_59_1334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3093_ net129 net24 _0842_ _0849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_71_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ _0494_ clknet_leaf_64_core_clock dmmu1.page_table\[4\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6189__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6852_ _0425_ clknet_leaf_33_core_clock dmmu0.page_table\[1\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5803_ _2806_ _0406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4739__A2 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ _0356_ clknet_leaf_41_core_clock dmmu1.page_table\[13\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3995_ _1655_ _1656_ _1439_ _1657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5734_ _2057_ _2760_ _2762_ net980 _2764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5665_ _2723_ _0351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4616_ _2098_ _0736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5164__A2 _2429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5596_ _2451_ _2681_ _2684_ net851 _2686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4547_ _2056_ _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4911__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3464__I _1203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input261_I dcache_wb_o_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input359_I ic1_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6113__A1 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4478_ _2012_ _0684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6217_ _0599_ clknet_leaf_83_core_clock immu_1.page_table\[7\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3429_ _1154_ _1169_ _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_22_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5872__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6148_ _3004_ _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_13_Left_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6079_ _2786_ _2958_ _2960_ net989 _2964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4427__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5624__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4978__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3650__A2 net242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5927__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6601__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_2049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output480_I net480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5155__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6751__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3307__C _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4666__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4418__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5091__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3641__A2 net262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3549__I _1274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6281__CLK clknet_leaf_36_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5394__A2 _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3780_ immu_1.page_table\[10\]\[1\] immu_1.page_table\[11\]\[1\] _1404_ _1449_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5450_ _1891_ _1892_ _2599_ _2600_ _2601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_2_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4401_ _1858_ _1957_ _1959_ net777 _1965_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_2034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput504 net504 c1_i_req_data[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5381_ _2561_ _0229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput515 net515 c1_i_req_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput526 net526 dcache_mem_addr[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput537 net537 dcache_mem_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7120_ net59 net582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput548 net548 dcache_mem_i_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4332_ _1924_ _0626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput559 net559 dcache_mem_req vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7051_ net287 net438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_49_core_clock clknet_3_6_0_core_clock clknet_leaf_49_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4263_ _1855_ _1876_ _1878_ net850 _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6002_ _2919_ _0492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3214_ dmmu1.page_table\[0\]\[2\] dmmu1.page_table\[1\]\[2\] dmmu1.page_table\[2\]\[2\]
+ dmmu1.page_table\[3\]\[2\] _0899_ _0931_ _0962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_78_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4121__A3 _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4194_ _1826_ _1828_ _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3145_ net106 net158 _0894_ _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__4409__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5606__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3076_ net220 _0831_ _0839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6624__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6904_ _0477_ clknet_leaf_59_core_clock dmmu1.page_table\[5\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input107_I c1_o_c_instr_long vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6835_ _0408_ clknet_leaf_46_core_clock dmmu1.page_table\[9\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5909__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6766_ _0339_ clknet_leaf_31_core_clock dmmu0.page_table\[5\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_1769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3978_ _1375_ _1640_ _1641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6774__CLK clknet_leaf_102_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3396__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4593__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5717_ _2753_ _0373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6697_ _0270_ clknet_leaf_32_core_clock dmmu0.page_table\[4\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5137__A2 _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5648_ net95 _2698_ _2700_ net788 _2714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_88_core_clock clknet_3_4_0_core_clock clknet_leaf_88_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6185__I1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input72_I c0_o_req_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5579_ _2101_ _2664_ _2666_ net1044 _2675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4896__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold240 dmmu0.page_table\[9\]\[7\] net974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold251 immu_1.page_table\[6\]\[7\] net985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold262 dmmu1.page_table\[14\]\[11\] net996 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold273 immu_1.page_table\[14\]\[7\] net1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold284 dmmu1.page_table\[0\]\[11\] net1018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold295 immu_1.page_table\[2\]\[8\] net1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4648__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_2298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4820__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3623__A2 net268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5376__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3482__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5128__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3234__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6089__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5836__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3311__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6647__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_2038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput8 c0_o_instr_long_addr[3] net8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_1296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4950_ _2269_ _2299_ _2302_ dmmu0.page_table\[7\]\[3\] _2306_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_1602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3901_ _1564_ _1565_ _1367_ _1566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6797__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4881_ _2256_ _0034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6013__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6620_ _0193_ clknet_leaf_15_core_clock immu_0.page_table\[0\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3832_ immu_1.page_table\[4\]\[3\] immu_1.page_table\[5\]\[3\] immu_1.page_table\[6\]\[3\]
+ immu_1.page_table\[7\]\[3\] _1435_ _1469_ _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_6_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3378__A1 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6551_ _0124_ clknet_leaf_20_core_clock immu_0.page_table\[6\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3763_ _1375_ _1428_ _1431_ _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_12_1977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5502_ _2631_ _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3473__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6482_ _0055_ clknet_leaf_28_core_clock dmmu0.page_table\[7\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3694_ _1337_ net233 _1365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4327__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5433_ _2591_ _0251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3225__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4878__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5364_ _1996_ _2535_ _2537_ dmmu0.page_table\[15\]\[12\] _2551_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7103_ net211 net563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4315_ _1846_ _1911_ _1914_ immu_1.page_table\[2\]\[1\] _1916_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5295_ _1814_ _2502_ _2504_ immu_0.page_table\[0\]\[7\] _2511_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_22_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7034_ net299 net450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4246_ _1870_ _1840_ _1842_ immu_1.page_table\[9\]\[10\] _1871_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4177_ _1815_ _1792_ _1794_ net988 _1816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input224_I dcache_mem_o_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3128_ net18 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_2_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5669__I _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3059_ net227 _0822_ _0830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4802__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3161__S0 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3189__I _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _0391_ clknet_leaf_67_core_clock dmmu1.page_table\[11\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5358__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6749_ _0322_ clknet_leaf_32_core_clock dmmu0.page_table\[6\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_2474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_2485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_2496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output443_I net443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7124__I net69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5818__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4097__A2 net383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3844__A2 net705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1078 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_38_Left_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_1343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3099__I _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_Left_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5521__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4100_ _1755_ _1756_ _1757_ net704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5080_ _2380_ _0109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_36_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_10_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5285__A1 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4031_ _1416_ _1691_ _1692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_1860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5037__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_56_Left_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5982_ _2908_ _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3599__A1 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4933_ _1796_ _2285_ _2287_ _1845_ _2293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4864_ _1803_ _2242_ _2244_ dmmu0.page_table\[9\]\[3\] _2248_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_13 net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_24 _1268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3815_ _0813_ _1482_ _1483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6603_ _0176_ clknet_leaf_5_core_clock immu_0.page_table\[1\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4795_ _2154_ _2205_ _2206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_43_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6534_ _0107_ clknet_leaf_2_core_clock immu_0.page_table\[8\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ net368 _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_6_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_65_Left_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6465_ _0038_ clknet_leaf_22_core_clock dmmu0.page_table\[8\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3677_ _1337_ net252 _1352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6812__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input174_I c1_o_req_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5416_ _1977_ _2468_ _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6396_ _0778_ clknet_leaf_104_core_clock immu_0.page_table\[15\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5347_ _2542_ _0214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4720__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input341_I ic1_mem_data[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5278_ _1789_ _1973_ _2501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6962__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input35_I c0_o_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4229_ _1858_ _1841_ _1843_ net876 _1859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_74_Left_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_1906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_2028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4251__A2 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_2039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6342__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_inner_730 c1_i_core_int_sreg[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7119__I net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5200__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3762__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6492__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5503__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_1_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5267__A1 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3373__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5019__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_76_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Left_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4778__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_48_1661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4941__I _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3557__I _1278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3600_ _1300_ net427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput11 c0_o_instr_long_addr[6] net11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput22 c0_o_mem_addr[3] net22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4580_ _2078_ _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5742__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput33 c0_o_mem_data[13] net33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_80_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput44 c0_o_mem_data[9] net44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3531_ net143 net38 _0850_ _1265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput55 c0_o_mem_sel[0] net55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4950__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput66 c0_o_req_addr[1] net66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput77 c0_sr_bus_addr[10] net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_57_1908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput88 c0_sr_bus_addr[6] net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6250_ _0632_ clknet_leaf_83_core_clock immu_1.page_table\[5\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput99 c0_sr_bus_data_o[4] net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3462_ _0894_ _1191_ _1192_ _0895_ _1201_ _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_58_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6985__CLK clknet_leaf_73_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3505__A1 _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5201_ _2454_ _0156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4702__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6181_ dmmu1.long_off_reg\[5\] _1858_ _3016_ _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_1280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3393_ _0906_ _1134_ _1135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5132_ _2332_ _2397_ _2399_ net758 _2411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_4_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6215__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5063_ _2267_ _2367_ _2369_ immu_0.page_table\[8\]\[2\] _2372_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4014_ _1366_ _1675_ _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3241__B _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6365__CLK clknet_leaf_75_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5965_ _2792_ _2890_ _2892_ dmmu1.page_table\[5\]\[6\] _2899_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3036__A3 _0815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5430__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4916_ _2280_ _0045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5896_ _2860_ _0445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5981__A2 _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4847_ _1821_ _2223_ _2225_ net792 _2237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3419__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input291_I ic0_mem_data[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input389_I inner_wb_i_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5194__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4778_ _1803_ _2191_ _2193_ immu_0.page_table\[12\]\[3\] _2197_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6517_ _0090_ clknet_leaf_0_core_clock immu_0.page_table\[9\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3729_ _1394_ _1395_ _1398_ _1372_ _1366_ _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_TAPCELL_ROW_73_2400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_73_2411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6448_ _0021_ clknet_leaf_10_core_clock dmmu0.page_table\[10\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5497__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6379_ _0761_ clknet_leaf_74_core_clock immu_1.page_table\[11\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput404 inner_wb_i_dat[9] net404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_25_1998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_2204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6708__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_2226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output406_I net406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6858__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3983__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6238__CLK clknet_leaf_91_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6388__CLK clknet_leaf_72_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3346__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4463__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3266__A3 _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ _2103_ _2760_ _2762_ dmmu1.page_table\[11\]\[9\] _2772_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_1413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5963__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4701_ _2149_ _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5681_ _2733_ _0357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4632_ _1912_ _2107_ _2109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5176__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4074__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4563_ _1860_ _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_29_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6302_ _0684_ clknet_leaf_93_core_clock immu_1.page_table\[1\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3514_ dmmu1.page_table\[4\]\[12\] dmmu1.page_table\[5\]\[12\] dmmu1.page_table\[6\]\[12\]
+ dmmu1.page_table\[7\]\[12\] _0886_ _0900_ _1252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_40_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4494_ _2022_ _0690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5479__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6233_ _0615_ clknet_leaf_81_core_clock immu_1.page_table\[0\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3445_ _1180_ _1183_ _1184_ _1185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6164_ _3012_ _0561_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3376_ _0879_ _1112_ _1117_ _0860_ _1118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_5115_ _2402_ _0122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6095_ net199 _2957_ _2959_ net924 _2972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input137_I c1_o_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5046_ _2361_ _0094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input304_I ic0_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6997_ _0570_ clknet_leaf_95_core_clock dmmu1.long_off_reg\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_24_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5948_ _2888_ _0469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3965__A1 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ net209 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_62_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4509__A3 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5706__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4142__A1 net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput201 c1_sr_bus_data_o[1] net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6530__CLK clknet_leaf_1_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput212 dcache_mem_ack net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_output523_I net523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput223 dcache_mem_o_data[3] net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput234 dcache_wb_adr[12] net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_1659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput245 dcache_wb_adr[22] net245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7132__I net62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput256 dcache_wb_o_dat[0] net256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput267 dcache_wb_o_dat[5] net267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3328__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput278 ic0_mem_data[10] net278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput289 ic0_mem_data[20] net289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4445__A2 _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5642__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6680__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5945__A2 _2872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3500__S0 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4056__S1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4905__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3835__I _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3803__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4381__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_39_core_clock clknet_3_6_0_core_clock clknet_leaf_39_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3230_ _0975_ _0976_ _0938_ _0977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3161_ dmmu1.page_table\[0\]\[0\] dmmu1.page_table\[1\]\[0\] dmmu1.page_table\[2\]\[0\]
+ dmmu1.page_table\[3\]\[0\] _0908_ _0910_ _0911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__7042__I net278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3092_ _0848_ net536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6920_ _0493_ clknet_leaf_63_core_clock dmmu1.page_table\[4\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6851_ _0424_ clknet_leaf_36_core_clock dmmu0.page_table\[1\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _2782_ _2802_ _2804_ net960 _2806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3994_ immu_1.page_table\[0\]\[8\] immu_1.page_table\[1\]\[8\] immu_1.page_table\[2\]\[8\]
+ immu_1.page_table\[3\]\[8\] _1404_ _1540_ _1656_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6782_ _0355_ clknet_leaf_45_core_clock dmmu1.page_table\[13\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3947__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ _2763_ _0379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6403__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5149__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5664_ dmmu0.long_off_reg\[6\] _1812_ _2716_ _2723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_78_core_clock clknet_3_5_0_core_clock clknet_leaf_78_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4615_ _2065_ _2090_ _2092_ net809 _2098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5595_ _2685_ _0319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3745__I net369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4546_ _2051_ _2053_ _2055_ net871 _2056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6553__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4477_ net198 _1998_ _2000_ immu_1.page_table\[1\]\[10\] _2012_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_40_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6113__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input254_I dcache_wb_adr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4124__A1 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5321__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6216_ _0598_ clknet_leaf_89_core_clock immu_1.page_table\[7\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3428_ _1159_ _1168_ _0821_ _1169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5872__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6147_ _1845_ _3000_ _3002_ net817 _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3480__I _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3359_ _0938_ _1101_ _0958_ _1102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6078_ _2963_ _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5624__A1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4427__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5029_ _1790_ _2240_ _2351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5927__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7127__I net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4363__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output640_I net640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4666__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_15_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6426__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3929__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6576__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7037__I net304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4400_ _1964_ _0654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3788__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5551__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5380_ _2459_ _2553_ _2555_ dmmu0.page_table\[11\]\[5\] _2561_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput505 net505 c1_i_req_data[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput516 net516 c1_i_req_data_valid vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput527 net527 dcache_mem_addr[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_50_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4331_ _1868_ _1911_ _1914_ immu_1.page_table\[2\]\[9\] _1924_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput538 net538 dcache_mem_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput549 net549 dcache_mem_i_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5780__I _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7050_ net286 net437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4106__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4262_ _1882_ _0598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6001_ _2849_ _2907_ _2909_ dmmu1.page_table\[4\]\[9\] _2919_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3213_ _0959_ _0960_ _0884_ _0961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_78_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4193_ _1827_ net181 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3144_ net158 _0893_ _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_39_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3960__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4409__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5606__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5457__I1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3075_ _0838_ net472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_1018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ _0476_ clknet_leaf_53_core_clock dmmu1.page_table\[5\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6834_ _0407_ clknet_leaf_47_core_clock dmmu1.page_table\[9\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5909__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6031__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6919__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6765_ _0338_ clknet_leaf_13_core_clock dmmu0.page_table\[5\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3977_ immu_0.page_table\[12\]\[7\] immu_0.page_table\[13\]\[7\] immu_0.page_table\[14\]\[7\]
+ immu_0.page_table\[15\]\[7\] _1487_ _1390_ _1640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4593__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3396__A2 _1128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5716_ _2069_ _2743_ _2745_ net1068 _2753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6696_ _0269_ clknet_leaf_31_core_clock dmmu0.page_table\[4\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5647_ _2713_ _0343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input371_I ic1_wb_adr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3779__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5578_ _2674_ _0313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input65_I c0_o_req_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold230 immu_1.page_table\[4\]\[8\] net964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4896__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold241 dmmu1.page_table\[12\]\[10\] net975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4529_ _1866_ _2033_ _2035_ dmmu1.page_table\[14\]\[8\] _2044_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold252 dmmu1.page_table\[1\]\[6\] net986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold263 dmmu0.page_table\[4\]\[3\] net997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold274 immu_0.page_table\[10\]\[10\] net1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold285 dmmu0.page_table\[1\]\[0\] net1019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold296 dmmu1.page_table\[11\]\[4\] net1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_6_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_2299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7179_ net398 net651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_1776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_6_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3871__A3 _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6449__CLK clknet_leaf_99_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5073__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3703__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_2073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6599__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5781__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3318__C _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6089__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_2090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5836__A1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3311__A2 _1055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 c0_o_instr_long_addr[4] net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3900_ _1384_ immu_0.page_table\[12\]\[5\] _1390_ _1565_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_1636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4880_ _1994_ _2241_ _2243_ dmmu0.page_table\[9\]\[11\] _2256_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_54_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6013__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3831_ _1368_ _1491_ _1497_ _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_12_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4575__A1 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3762_ _1372_ _1381_ _1430_ _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6550_ _0123_ clknet_leaf_3_core_clock immu_0.page_table\[6\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5772__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5501_ _2300_ _2629_ _2631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_70_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6481_ _0054_ clknet_leaf_29_core_clock dmmu0.page_table\[7\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3693_ _1350_ net311 _1360_ _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_1680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4327__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5432_ _2461_ _2582_ _2584_ net855 _2591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_83_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4878__A2 _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5363_ _2550_ _0222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7102_ net211 net517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4314_ _1915_ _0617_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_1175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5294_ _2510_ _0193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7033_ net288 net439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4245_ net198 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4176_ _1814_ _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3933__S0 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3127_ _0876_ _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_2_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input217_I dcache_mem_o_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3066__A1 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3058_ _0829_ net479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6741__CLK clknet_leaf_42_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4263__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4802__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3161__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6817_ _0390_ clknet_leaf_42_core_clock dmmu1.page_table\[11\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_2092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6891__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6748_ _0321_ clknet_leaf_31_core_clock dmmu0.page_table\[6\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5763__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6679_ _0252_ clknet_leaf_33_core_clock dmmu0.page_table\[2\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5515__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_2475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_2497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5818__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output436_I net436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6271__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3924__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output603_I net603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7140__I net389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_2072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3057__A1 net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_1972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6614__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_55_1847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4030_ immu_1.page_table\[12\]\[9\] immu_1.page_table\[13\]\[9\] immu_1.page_table\[14\]\[9\]
+ immu_1.page_table\[15\]\[9\] _1409_ _1410_ _1691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5285__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Right_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6764__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4493__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7050__I net286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5037__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5981_ _1770_ _2906_ _2908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4932_ _2289_ _2292_ _1771_ _0049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3599__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5993__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4863_ _2247_ _0025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6602_ _0175_ clknet_leaf_6_core_clock immu_0.page_table\[2\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_14 net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_25 _1268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3814_ _1434_ net705 _1476_ _1481_ _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_12_1753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4794_ _2171_ net76 _2205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_27_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6533_ _0106_ clknet_leaf_0_core_clock immu_0.page_table\[8\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3745_ net369 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_15_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6464_ _0037_ clknet_leaf_23_core_clock dmmu0.page_table\[8\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3676_ _1350_ net322 _1326_ _1351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5415_ _2580_ _0244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6294__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6395_ _0777_ clknet_leaf_106_core_clock immu_0.page_table\[15\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4720__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input167_I c1_o_req_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5346_ _2455_ _2536_ _2538_ net1075 _2542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_71_2350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5277_ _1776_ _2500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input334_I ic1_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4228_ _1857_ _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_39_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3287__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input28_I c0_o_mem_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4159_ net98 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_58_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_2290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_2154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_2165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4251__A3 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4539__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_inner_720 c1_i_core_int_sreg[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_19_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_inner_731 c1_i_core_int_sreg[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_46_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5200__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_2537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6637__CLK clknet_leaf_10_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3762__A2 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6161__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7135__I net65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_1700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5267__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3278__A1 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4475__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3373__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3104__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5019__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4778__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 c0_o_instr_long_addr[7] net12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput23 c0_o_mem_addr[4] net23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput34 c0_o_mem_data[14] net34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput45 c0_o_mem_high_addr[0] net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3530_ _1264_ net551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4950__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4950__B2 dmmu0.page_table\[7\]\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput56 c0_o_mem_sel[1] net56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_1595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput67 c0_o_req_addr[2] net67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput78 c0_sr_bus_addr[11] net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput89 c0_sr_bus_addr[7] net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3461_ _0912_ _1195_ _1200_ _1201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7045__I net281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5200_ _2453_ _2447_ _2449_ net1003 _2454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4702__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6180_ _3021_ _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_1893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3392_ dmmu1.page_table\[8\]\[8\] dmmu1.page_table\[9\]\[8\] dmmu1.page_table\[10\]\[8\]
+ dmmu1.page_table\[11\]\[8\] _0887_ _0909_ _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_58_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5131_ _2410_ _0130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5062_ _2371_ _0100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3269__A1 net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4013_ immu_0.page_table\[12\]\[8\] immu_0.page_table\[13\]\[8\] immu_0.page_table\[14\]\[8\]
+ immu_0.page_table\[15\]\[8\] _1487_ _1390_ _1675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_79_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5964_ _2898_ _0475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5430__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4915_ _1819_ _2261_ _2263_ dmmu0.page_table\[8\]\[9\] _2280_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3441__A1 net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5895_ _2782_ _2856_ _2858_ net1081 _2860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5718__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4846_ _2236_ _0019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5194__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4777_ _2196_ _0799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input284_I ic0_mem_data[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6516_ _0089_ clknet_leaf_7_core_clock immu_0.page_table\[9\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3728_ _1385_ immu_0.page_table\[5\]\[0\] _1397_ _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_70_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6447_ _0020_ clknet_leaf_9_core_clock dmmu0.page_table\[10\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3659_ _1337_ net248 _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5497__A2 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6378_ _0760_ clknet_leaf_76_core_clock immu_1.page_table\[11\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5329_ net93 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5404__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4457__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_2205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_2216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_2105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4209__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3680__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5957__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_2086 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3983__A2 _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_29_core_clock clknet_3_3_0_core_clock clknet_leaf_29_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_37_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4696__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4999__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3346__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3671__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6802__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3423__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4700_ _2067_ _2139_ _2142_ net863 _2149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_57_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5680_ _2063_ _2726_ _2728_ dmmu1.page_table\[13\]\[4\] _2733_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6952__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4631_ _2107_ _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_leaf_68_core_clock clknet_3_6_0_core_clock clknet_leaf_68_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5176__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5783__I _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_22_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4562_ _2066_ _0714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ _0683_ clknet_leaf_81_core_clock immu_1.page_table\[1\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3513_ dmmu1.page_table\[0\]\[12\] dmmu1.page_table\[1\]\[12\] dmmu1.page_table\[2\]\[12\]
+ dmmu1.page_table\[3\]\[12\] _0886_ _0900_ _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_12_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4493_ _1858_ _2014_ _2016_ immu_1.page_table\[3\]\[5\] _2022_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5479__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6232_ _0614_ clknet_leaf_86_core_clock immu_1.page_table\[0\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3444_ _1180_ _1183_ _1119_ _1184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6163_ _2849_ _3000_ _3002_ net993 _3012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3375_ _1114_ _1116_ _0879_ _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5114_ _2265_ _2398_ _2400_ immu_0.page_table\[6\]\[1\] _2402_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6332__CLK clknet_leaf_75_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6094_ _2971_ _0532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4439__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5045_ _2275_ _2352_ _2354_ immu_0.page_table\[9\]\[6\] _2361_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3662__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6482__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5939__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6996_ _0569_ clknet_leaf_95_core_clock dmmu1.long_off_reg\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3414__A1 net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5947_ _2049_ _2872_ _2874_ net1067 _2888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4611__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5878_ _2848_ _0439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input95_I c0_sr_bus_data_o[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4829_ _1797_ _2224_ _2226_ dmmu0.page_table\[10\]\[1\] _2228_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3717__A2 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3427__B _1167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4678__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput202 c1_sr_bus_data_o[2] net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput213 dcache_mem_exception net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_21_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput224 dcache_mem_o_data[4] net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput235 dcache_wb_adr[13] net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput246 dcache_wb_adr[23] net246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput257 dcache_wb_o_dat[10] net257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput268 dcache_wb_o_dat[6] net268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output516_I net516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3328__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput279 ic0_mem_data[11] net279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6825__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5642__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3653__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6975__CLK clknet_leaf_102_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3500__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6205__CLK clknet_leaf_93_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4905__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6107__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4381__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6355__CLK clknet_leaf_71_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_88_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4133__A2 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5330__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3160_ _0909_ _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_20_1137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3892__A1 net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold1 ic0_wb_cyc net735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_55_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3091_ net128 net23 _0842_ _0848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4841__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _0423_ clknet_leaf_13_core_clock dmmu0.page_table\[1\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5801_ _2805_ _0405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5397__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6781_ _0354_ clknet_leaf_44_core_clock dmmu1.page_table\[13\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_8_Right_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3993_ immu_1.page_table\[4\]\[8\] immu_1.page_table\[5\]\[8\] immu_1.page_table\[6\]\[8\]
+ immu_1.page_table\[7\]\[8\] _1404_ _1540_ _1655_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5732_ _2051_ _2760_ _2762_ dmmu1.page_table\[11\]\[0\] _2763_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3947__A2 _1594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_2019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5149__A1 _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5663_ _2722_ _0350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ _2097_ _0735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5594_ _2444_ _2681_ _2684_ dmmu0.page_table\[6\]\[0\] _2685_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4545_ _2054_ _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_40_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_2041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4476_ _2011_ _0683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6215_ _0597_ clknet_leaf_88_core_clock immu_1.page_table\[7\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4857__I _2243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5321__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4124__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3427_ _0912_ _1162_ _1167_ _0895_ _1168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XPHY_EDGE_ROW_39_Right_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_1936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6848__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input247_I dcache_wb_adr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5872__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6146_ _3003_ _0552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3358_ dmmu0.page_table\[8\]\[7\] dmmu0.page_table\[9\]\[7\] dmmu0.page_table\[10\]\[7\]
+ dmmu0.page_table\[11\]\[7\] _0950_ _0952_ _1101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__3883__A1 net111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6077_ _2784_ _2958_ _2960_ net912 _2963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3289_ dmmu0.page_table\[13\]\[4\] _1035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5085__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5624__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5028_ _2350_ _0087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3635__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input10_I c0_o_instr_long_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6998__CLK clknet_leaf_95_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_90_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6979_ _0552_ clknet_leaf_79_core_clock immu_1.page_table\[8\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_48_Right_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6228__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4060__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6378__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4899__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Right_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output633_I net633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7143__I net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_66_Right_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3485__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5551__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_75_Right_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3788__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_2096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput506 net506 c1_i_req_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput517 net517 c1_rst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput528 net528 dcache_mem_addr[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4330_ _1923_ _0625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput539 net539 dcache_mem_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4106__A2 net327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ _1852_ _1876_ _1878_ net769 _1882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6000_ _2918_ _0491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5854__A2 _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3212_ _0940_ _0883_ _0960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4192_ net188 _1827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input2_I c0_o_c_instr_long vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3865__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3143_ net124 _0892_ _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3960__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5067__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5606__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3074_ net219 _0831_ _0838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3617__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4814__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _0475_ clknet_leaf_54_core_clock dmmu1.page_table\[5\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6833_ _0406_ clknet_leaf_48_core_clock dmmu1.page_table\[9\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3957__S _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6764_ _0337_ clknet_leaf_30_core_clock dmmu0.page_table\[5\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3976_ _1637_ _1638_ _1366_ _1639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6520__CLK clknet_leaf_109_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5715_ _2752_ _0372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4593__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5790__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _0268_ clknet_leaf_32_core_clock dmmu0.page_table\[4\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input197_I c1_sr_bus_data_o[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5646_ net94 _2698_ _2700_ dmmu0.page_table\[5\]\[11\] _2713_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3228__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4345__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3779__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5577_ _2069_ _2664_ _2666_ dmmu1.page_table\[15\]\[7\] _2674_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold220 immu_0.page_table\[3\]\[8\] net954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input364_I ic1_wb_adr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4528_ _2043_ _0703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold231 dmmu0.page_table\[10\]\[11\] net965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold242 immu_0.page_table\[14\]\[6\] net976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold253 dmmu1.page_table\[12\]\[0\] net987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input58_I c0_o_req_active vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold264 dmmu0.page_table\[3\]\[9\] net998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold275 immu_1.page_table\[6\]\[8\] net1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4459_ _1845_ _1999_ _2001_ immu_1.page_table\[1\]\[1\] _2003_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xhold286 immu_1.page_table\[9\]\[7\] net1020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold297 immu_0.page_table\[9\]\[4\] net1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7178_ net397 net650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3856__A1 net110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6129_ net213 net212 _2991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5412__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3608__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3703__S1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5211__I _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4033__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5230__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output583_I net583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5781__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3219__S0 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5533__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6089__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5297__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5836__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5049__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6543__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6013__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3830_ _1378_ _1381_ _1496_ _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_32_2073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4024__A1 net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3458__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5772__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3761_ _1368_ _1429_ _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4575__A2 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7048__I net284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6693__CLK clknet_leaf_89_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5500_ _2629_ _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_3_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ _0053_ clknet_leaf_30_core_clock dmmu0.page_table\[7\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3692_ _1348_ net365 _1363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5431_ _2590_ _0250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4327__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5362_ _1994_ _2535_ _2537_ net830 _2550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7101_ net330 net516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_80_1657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4313_ _1824_ _1911_ _1914_ immu_1.page_table\[2\]\[0\] _1915_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5293_ _1811_ _2502_ _2504_ immu_0.page_table\[0\]\[6\] _2510_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_26_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4200__I net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7032_ net277 net428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4244_ _1869_ _0593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3838__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4175_ net102 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3933__S1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3126_ _0875_ _0876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_2_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3260__B _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3057_ net226 _0822_ _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4263__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3066__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input112_I c1_o_instr_long_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_1174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6816_ _0389_ clknet_leaf_40_core_clock dmmu1.page_table\[11\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4015__A1 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5763__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6747_ _0320_ clknet_leaf_32_core_clock dmmu0.page_table\[6\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3959_ _1434_ _1621_ _1622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_1456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6678_ _0251_ clknet_leaf_35_core_clock dmmu0.page_table\[2\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5629_ _2704_ _0334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5515__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_2476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_2498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6416__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5818__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3829__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output429_I net429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3924__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6566__CLK clknet_leaf_18_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3057__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_2079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5876__I net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5203__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5754__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3860__S0 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_27_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4493__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5690__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3540__I0 net147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5980_ _2906_ _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5442__B1 _2583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ _1776_ _2290_ _2291_ _1823_ _2292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5993__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4862_ _1800_ _2242_ _2244_ net773 _2247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6601_ _0174_ clknet_leaf_16_core_clock immu_0.page_table\[2\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3813_ _1433_ _1477_ _1480_ _1415_ _1481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA_15 net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _2204_ _0807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6532_ _0105_ clknet_leaf_1_core_clock immu_0.page_table\[8\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3744_ immu_1.page_table\[12\]\[0\] immu_1.page_table\[13\]\[0\] immu_1.page_table\[14\]\[0\]
+ immu_1.page_table\[15\]\[0\] _1409_ _1410_ _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_12_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _0036_ clknet_leaf_27_core_clock dmmu0.page_table\[8\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3675_ _0813_ _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_42_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6439__CLK clknet_leaf_21_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5414_ immu_0.high_addr_off\[7\] _1815_ _2572_ _2580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6394_ _0776_ clknet_leaf_105_core_clock immu_0.page_table\[15\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5345_ _2541_ _0213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4720__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_2340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5276_ _2499_ _0186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6589__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4227_ net205 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3531__I0 net143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input327_I ic0_wb_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ _1801_ _0575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_69_2280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3109_ net19 _0858_ _0859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_69_2291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4089_ net116 immu_1.high_addr_off\[6\] _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_2144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_2077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4539__A2 _2032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5736__B2 dmmu1.page_table\[11\]\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_inner_710 c0_i_core_int_sreg[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_inner_721 c1_i_core_int_sreg[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_inner_732 c1_i_core_int_sreg[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_30_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_19_core_clock clknet_3_2_0_core_clock clknet_leaf_19_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6161__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7151__I net391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4475__A1 net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5672__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5424__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4778__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A1 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_58_core_clock clknet_3_7_0_core_clock clknet_leaf_58_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput13 c0_o_mem_addr[0] net13 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3833__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput24 c0_o_mem_addr[5] net24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput35 c0_o_mem_data[15] net35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_1763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput46 c0_o_mem_high_addr[1] net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_80_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4950__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput57 c0_o_mem_we net57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput68 c0_o_req_addr[3] net68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput79 c0_sr_bus_addr[12] net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3460_ net123 _1197_ _1199_ _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_64_1449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6731__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4702__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3790__S _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3391_ _0896_ _1132_ _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5130_ _2330_ _2398_ _2400_ immu_0.page_table\[6\]\[9\] _2410_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_1758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4685__I _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5061_ _2265_ _2367_ _2369_ immu_0.page_table\[8\]\[1\] _2371_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6881__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4012_ _1367_ _1673_ _1674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_97_core_clock clknet_3_1_0_core_clock clknet_leaf_97_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5963_ _2790_ _2890_ _2892_ dmmu1.page_table\[5\]\[5\] _2898_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4914_ _2279_ _0044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5894_ _2859_ _0444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_95_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4845_ _1819_ _2224_ _2226_ dmmu0.page_table\[10\]\[9\] _2236_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5718__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6261__CLK clknet_leaf_83_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4776_ _1800_ _2191_ _2193_ immu_0.page_table\[12\]\[2\] _2196_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5194__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3824__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6515_ _0088_ clknet_leaf_8_core_clock immu_0.page_table\[9\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3727_ _1396_ immu_0.page_table\[4\]\[0\] _1397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_47_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3764__I _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input277_I ic0_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6143__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6446_ _0019_ clknet_leaf_12_core_clock dmmu0.page_table\[10\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3658_ inner_wb_arbiter.o_sel_sig _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_30_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6377_ _0759_ clknet_leaf_73_core_clock immu_1.page_table\[11\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3589_ net216 _1219_ _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_64_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5328_ _2530_ _0207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input40_I c0_o_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5259_ _1799_ _2486_ _2488_ immu_0.page_table\[1\]\[2\] _2491_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4457__A1 _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4209__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3680__A2 net323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6604__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output496_I net496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3196__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output663_I net663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7146__I net401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4696__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5893__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4448__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4999__A2 _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A2 net251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6284__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3785__S _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4059__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4630_ _1838_ _1892_ _2028_ _2107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5176__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4561_ _2065_ _2053_ _2055_ net826 _2066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _0682_ clknet_leaf_86_core_clock immu_1.page_table\[1\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3512_ net157 dmmu1.long_off_reg\[7\] _1249_ _1250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_44_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6125__A1 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4492_ _2021_ _0689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6231_ _0613_ clknet_leaf_83_core_clock immu_1.page_table\[0\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3443_ _1142_ _1181_ _1182_ _1183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_29_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6162_ _3011_ _0560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3374_ _0940_ _1115_ _1116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5113_ _2401_ _0121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6093_ _2851_ _2957_ _2959_ dmmu1.page_table\[1\]\[10\] _2971_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5304__I _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4439__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5636__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5044_ _2360_ _0093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3252__C _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3111__A1 net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6627__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3662__A2 net319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5939__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6995_ _0568_ clknet_leaf_95_core_clock dmmu1.long_off_reg\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6061__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5946_ _2887_ _0468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4611__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6777__CLK clknet_leaf_100_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5877_ _2847_ _2836_ _2838_ dmmu1.page_table\[8\]\[8\] _2848_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input394_I inner_wb_i_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4828_ _2227_ _0010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4375__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input88_I c0_sr_bus_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4759_ _1815_ _2175_ _2177_ net1076 _2185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3427__C _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6429_ _0002_ clknet_leaf_104_core_clock immu_0.page_table\[13\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4678__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3350__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput203 c1_sr_bus_data_o[3] net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput214 dcache_mem_o_data[0] net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xinput225 dcache_mem_o_data[5] net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5214__I _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput236 dcache_wb_adr[14] net236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput247 dcache_wb_adr[2] net247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput258 dcache_wb_o_dat[11] net258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput269 dcache_wb_o_dat[7] net269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output509_I net509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3653__A2 net317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_core_clock clknet_3_1_0_core_clock clknet_leaf_9_core_clock vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_54_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3169__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4905__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6107__A1 _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5866__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5330__A2 _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_105_core_clock clknet_3_0_0_core_clock clknet_leaf_105_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold2 icore_sregs.c1_disable net736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3090_ _0847_ net535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4841__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6043__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5800_ _2776_ _2802_ _2804_ net764 _2805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6780_ _0353_ clknet_leaf_45_core_clock dmmu1.page_table\[13\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3992_ _1651_ _1652_ _1653_ _1654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5397__A2 net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5731_ _2761_ _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5662_ dmmu0.long_off_reg\[5\] _1809_ _2716_ _2722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5149__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4357__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4613_ _2063_ _2090_ _2092_ immu_1.page_table\[13\]\[4\] _2097_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5593_ _2683_ _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_4_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4544_ _1912_ _2052_ _2054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3247__C _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4475_ net209 _1999_ _2001_ immu_1.page_table\[1\]\[9\] _2011_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_42_2031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6214_ _0596_ clknet_leaf_84_core_clock immu_1.page_table\[7\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3426_ _1164_ _1166_ net123 _1167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__5321__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6145_ _1823_ _3000_ _3002_ net1012 _3003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3357_ _0940_ _1099_ _1100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input142_I c1_o_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6076_ _2962_ _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3288_ _0882_ _1032_ _1033_ _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5085__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5027_ _2332_ _2336_ _2338_ net1008 _2350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3635__A2 net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4094__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5388__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6978_ _0551_ clknet_leaf_103_core_clock mem_dcache_arb.transfer_active vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3238__I2 dmmu1.page_table\[14\]\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3399__A1 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5929_ _2786_ _2873_ _2875_ net790 _2879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4899__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3571__A1 net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output459_I net459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5848__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__I net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6942__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3901__B _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_2066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6025__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4587__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3929__A3 _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3485__S1 _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6179__I1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4339__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5551__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput507 net507 c1_i_req_data[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput518 net518 dcache_mem_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_10_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_2059 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput529 net529 dcache_mem_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6472__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4260_ _1881_ _0597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3211_ _0956_ _0957_ _0958_ _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4191_ net190 _1825_ _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_24_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3142_ _0890_ _0891_ _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5067__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_2013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3073_ _0837_ net471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4814__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3617__A2 net265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6901_ _0474_ clknet_leaf_50_core_clock dmmu1.page_table\[5\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3173__S0 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_34_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6832_ _0405_ clknet_leaf_47_core_clock dmmu1.page_table\[9\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6763_ _0336_ clknet_leaf_29_core_clock dmmu0.page_table\[5\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3975_ immu_0.page_table\[4\]\[7\] immu_0.page_table\[5\]\[7\] immu_0.page_table\[6\]\[7\]
+ immu_0.page_table\[7\]\[7\] _1396_ _1371_ _1638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_50_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5714_ _2067_ _2743_ _2745_ net909 _2752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6694_ _0267_ clknet_leaf_31_core_clock dmmu0.page_table\[4\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_17_Left_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5645_ _2712_ _0342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3228__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6815__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5576_ _2673_ _0312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold210 immu_1.page_table\[15\]\[6\] net944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold221 immu_0.page_table\[8\]\[7\] net955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4527_ _1864_ _2033_ _2035_ dmmu1.page_table\[14\]\[7\] _2043_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3772__I net366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold232 dmmu1.page_table\[0\]\[9\] net966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold243 dmmu1.page_table\[4\]\[6\] net977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold254 immu_0.page_table\[11\]\[7\] net988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold265 dmmu1.page_table\[5\]\[0\] net999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input357_I ic1_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4458_ _2002_ _0674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold276 immu_0.page_table\[2\]\[7\] net1010 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold287 immu_0.page_table\[2\]\[3\] net1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold298 immu_0.page_table\[14\]\[2\] net1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3305__A1 net150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3409_ dmmu0.page_table\[0\]\[9\] dmmu0.page_table\[1\]\[9\] dmmu0.page_table\[2\]\[9\]
+ dmmu0.page_table\[3\]\[9\] _0863_ _0866_ _1150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7177_ net396 net649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4389_ _1912_ _1956_ _1958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6128_ _2990_ _0547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6059_ _2847_ _2941_ _2943_ net984 _2952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3608__A2 net274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6345__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4569__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5230__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5781__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3219__S1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6495__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5533__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7154__I net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5297__A1 net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5049__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_1798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5221__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3458__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6838__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3083__I0 net118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3760_ immu_0.page_table\[2\]\[1\] immu_0.page_table\[3\]\[1\] immu_0.page_table\[10\]\[1\]
+ immu_0.page_table\[11\]\[1\] _1424_ _1377_ _1429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_54_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5772__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4575__A3 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3783__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4980__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3691_ _1359_ _1361_ _1362_ net661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3793__S _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5430_ _2459_ _2582_ _2584_ net968 _2590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6988__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4732__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5361_ _2549_ _0221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7100_ net355 net508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4312_ _1913_ _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_1767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5292_ _2509_ _0192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7031_ net406 net409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4243_ _1868_ _1841_ _1843_ net1089 _1869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4174_ _1813_ _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3125_ net17 _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_39_1516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6368__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3056_ _0828_ net478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4263__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input105_I c0_sr_bus_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6815_ _0388_ clknet_leaf_65_core_clock dmmu1.page_table\[11\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6746_ _0319_ clknet_leaf_30_core_clock dmmu0.page_table\[6\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5763__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3958_ immu_1.page_table\[12\]\[7\] immu_1.page_table\[13\]\[7\] immu_1.page_table\[14\]\[7\]
+ immu_1.page_table\[15\]\[7\] _1441_ _1442_ _1621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3889_ net6 immu_0.high_addr_off\[1\] _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6677_ _0250_ clknet_leaf_13_core_clock dmmu0.page_table\[2\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5628_ _1799_ _2699_ _2701_ net746 _2704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5515__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input70_I c0_o_req_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_2477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_2488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5559_ _1874_ _2028_ _2031_ _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_76_2499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_1108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5451__A1 _1834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3462__B1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5203__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_48_core_clock clknet_3_6_0_core_clock clknet_leaf_48_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_1182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7149__I net404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_2_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4962__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3860__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6510__CLK clknet_leaf_2_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4493__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5690__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3540__I1 net42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_87_core_clock clknet_3_4_0_core_clock clknet_leaf_87_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5442__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4971__I _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ _1829_ _1837_ _2286_ _2291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__6660__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5993__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _2246_ _0024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_25_Left_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6600_ _0173_ clknet_leaf_17_core_clock immu_0.page_table\[2\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3812_ _1433_ _1478_ _1479_ _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_7_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4792_ _1821_ _2190_ _2192_ immu_0.page_table\[12\]\[10\] _2204_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_27_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_16 net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3300__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3743_ immu_1.page_table\[4\]\[0\] immu_1.page_table\[5\]\[0\] immu_1.page_table\[6\]\[0\]
+ immu_1.page_table\[7\]\[0\] _1409_ _1410_ _1413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6531_ _0104_ clknet_leaf_109_core_clock immu_0.page_table\[8\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6462_ _0035_ clknet_leaf_99_core_clock dmmu0.page_table\[9\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3674_ _1348_ net376 _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5413_ _2579_ _0243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6393_ _0775_ clknet_leaf_106_core_clock immu_0.page_table\[15\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5344_ _2453_ _2536_ _2538_ dmmu0.page_table\[15\]\[2\] _2541_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_1444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_71_2341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_34_Left_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_71_2352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5275_ net93 _2485_ _2487_ immu_0.page_table\[1\]\[10\] _2499_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_23_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4226_ _1856_ _0588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5130__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3531__I1 net38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4157_ _1800_ _1792_ _1794_ net938 _1801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input222_I dcache_mem_o_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3119__S0 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3108_ _0856_ _0857_ _0858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_2270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4088_ _1350_ _1579_ _1746_ _1747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_69_2292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3039_ mem_dcache_arb.select _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_2156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_43_Left_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_2034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5197__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinterconnect_inner_711 c0_i_core_int_sreg[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_18_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinterconnect_inner_722 c1_i_core_int_sreg[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_inner_733 c1_i_core_int_sreg[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_22_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4944__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6729_ _0302_ clknet_leaf_37_core_clock dmmu0.page_table\[3\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_22_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6161__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Left_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_1773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6533__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output441_I net441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput690 net690 inner_wb_o_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3358__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3181__B _0929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5672__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4475__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6683__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5424__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Left_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_1244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A2 _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_29_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4935__B1 _2291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput14 c0_o_mem_addr[10] net14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3833__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput25 c0_o_mem_addr[6] net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput36 c0_o_mem_data[1] net36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput47 c0_o_mem_high_addr[2] net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_52_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput58 c0_o_req_active net58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_70_Left_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput69 c0_o_req_addr[4] net69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3390_ dmmu1.page_table\[12\]\[8\] dmmu1.page_table\[13\]\[8\] dmmu1.page_table\[14\]\[8\]
+ dmmu1.page_table\[15\]\[8\] _0887_ _0909_ _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_0_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3910__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5060_ _2370_ _0099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5112__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4011_ immu_0.page_table\[8\]\[8\] immu_0.page_table\[9\]\[8\] immu_0.page_table\[10\]\[8\]
+ immu_0.page_table\[11\]\[8\] _1487_ _1390_ _1673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_74_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5962_ _2897_ _0474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4913_ _1817_ _2261_ _2263_ dmmu0.page_table\[8\]\[8\] _2279_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5893_ _2776_ _2856_ _2858_ dmmu1.page_table\[7\]\[0\] _2859_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_60_2020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_16_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5718__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4844_ _2235_ _0018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3729__B2 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4775_ _2195_ _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3824__S1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6514_ _0087_ clknet_leaf_105_core_clock immu_0.page_table\[10\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3726_ _1369_ _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_31_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6556__CLK clknet_leaf_18_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_2403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6445_ _0018_ clknet_leaf_23_core_clock dmmu0.page_table\[10\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3657_ _0814_ net318 _1326_ _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_1940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input172_I c1_o_req_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3588_ _1294_ net412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6376_ _0758_ clknet_leaf_74_core_clock immu_1.page_table\[11\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5327_ _2529_ _2516_ _2518_ net783 _2530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5103__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5258_ _2490_ _0177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input33_I c0_o_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4457__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4209_ _1824_ _1841_ _1843_ immu_1.page_table\[9\]\[0\] _1844_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5189_ _1780_ _1971_ _2445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_67_2207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_2218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_2229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3760__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_2107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4209__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3221__S _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5500__I _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4116__I _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output489_I net489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4393__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5342__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_5_Left_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5893__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4696__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7162__I net176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4448__A2 _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6429__CLK clknet_leaf_104_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3959__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_39_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4059__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6579__CLK clknet_leaf_3_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4908__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4560_ _1857_ _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5581__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_1334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3511_ _1216_ _1247_ _1248_ _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4491_ _1855_ _2014_ _2016_ net867 _2021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6125__A2 _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3442_ net49 dmmu0.long_off_reg\[4\] _1182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6230_ _0612_ clknet_leaf_80_core_clock immu_1.page_table\[0\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3373_ dmmu0.page_table\[4\]\[8\] dmmu0.page_table\[5\]\[8\] dmmu0.page_table\[6\]\[8\]
+ dmmu0.page_table\[7\]\[8\] _0864_ _0941_ _1115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6161_ _2847_ _3000_ _3002_ immu_1.page_table\[8\]\[8\] _3011_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7072__I net356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5112_ _2258_ _2398_ _2400_ immu_0.page_table\[6\]\[0\] _2401_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6092_ _2970_ _0531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5636__A1 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4439__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5043_ _2273_ _2352_ _2354_ immu_0.page_table\[9\]\[5\] _2360_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3105__I _0855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3111__A2 net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3742__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_2039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6994_ _0567_ clknet_leaf_95_core_clock dmmu1.long_off_reg\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5939__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6061__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5945_ _2047_ _2872_ _2874_ net840 _2887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4611__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3976__S _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5876_ net208 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_36_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4827_ _1777_ _2224_ _2226_ dmmu0.page_table\[10\]\[0\] _2227_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_2094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input387_I inner_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4375__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4758_ _2184_ _0792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_1423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3709_ _1375_ _1376_ _1378_ _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4689_ _2143_ _0764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4127__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5324__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6428_ _0001_ clknet_leaf_106_core_clock immu_0.page_table\[13\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_41_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4678__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6359_ _0741_ clknet_leaf_70_core_clock immu_1.page_table\[13\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3216__S _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput204 c1_sr_bus_data_o[4] net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3350__A2 _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput215 dcache_mem_o_data[10] net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput226 dcache_mem_o_data[6] net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput237 dcache_wb_adr[15] net237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput248 dcache_wb_adr[3] net248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput259 dcache_wb_o_dat[12] net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_58_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6721__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7157__I net171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5402__I1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6871__CLK clknet_leaf_48_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6107__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5315__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5866__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5618__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold3 immu_1.page_table\[0\]\[0\] net737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_59_1349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4841__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6043__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3991_ _1651_ _1652_ net107 _1653_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5730_ _2682_ _2759_ _2761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_18_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5661_ _2721_ _0349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7067__I net407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4357__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4612_ _2096_ _0734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5592_ _2682_ _2680_ _2683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_60_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ _2052_ _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_48_1754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4109__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4474_ _2010_ _0682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6213_ _0595_ clknet_leaf_82_core_clock immu_1.page_table\[7\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3425_ _0906_ _1165_ _1166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3356_ dmmu0.page_table\[12\]\[7\] dmmu0.page_table\[13\]\[7\] dmmu0.page_table\[14\]\[7\]
+ dmmu0.page_table\[15\]\[7\] _0882_ _0948_ _1099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6144_ _3001_ _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6075_ _2782_ _2958_ _2960_ dmmu1.page_table\[1\]\[1\] _2962_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3287_ _0882_ dmmu0.page_table\[14\]\[4\] _0941_ _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5085__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input135_I c1_o_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5026_ _2349_ _0086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6744__CLK clknet_leaf_40_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4293__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_2101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input302_I ic0_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _0550_ clknet_leaf_103_core_clock mem_dcache_arb.req0_pending vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4045__B1 _1705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5928_ _2878_ _0459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6894__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5859_ _2837_ _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_35_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5545__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4899__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3571__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5848__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5225__I _2469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output521_I net521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3706__S0 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4823__A2 _2222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6025__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4587__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5784__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4339__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6617__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput508 net508 c1_i_req_data[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput519 net519 dcache_mem_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_10_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3210_ net18 _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__4511__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4190_ net189 _1825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_24_1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3141_ net151 net150 net153 net152 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_59_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5067__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3072_ net218 _0831_ _0837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_59_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4814__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6900_ _0473_ clknet_leaf_52_core_clock dmmu1.page_table\[5\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3173__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_2009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6831_ _0404_ clknet_leaf_68_core_clock dmmu1.page_table\[10\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5775__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6762_ _0335_ clknet_leaf_46_core_clock dmmu0.page_table\[5\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3974_ immu_0.page_table\[0\]\[7\] immu_0.page_table\[1\]\[7\] immu_0.page_table\[2\]\[7\]
+ immu_0.page_table\[3\]\[7\] _1396_ _1371_ _1637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_9_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5713_ _2751_ _0371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6693_ _0266_ clknet_leaf_89_core_clock immu_1.high_addr_off\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3258__C _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5527__B1 _2631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5644_ _2531_ _2698_ _2700_ net742 _2712_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6297__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5575_ _2067_ _2664_ _2666_ dmmu1.page_table\[15\]\[6\] _2673_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold200 immu_1.page_table\[6\]\[4\] net934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold211 immu_1.page_table\[8\]\[7\] net945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_14_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4526_ _2042_ _0702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold222 dmmu1.page_table\[5\]\[12\] net956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold233 immu_1.page_table\[12\]\[5\] net967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold244 immu_0.page_table\[8\]\[0\] net978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold255 dmmu1.page_table\[1\]\[3\] net989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold266 dmmu1.page_table\[8\]\[3\] net1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4457_ _1823_ _1999_ _2001_ immu_1.page_table\[1\]\[0\] _2002_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xhold277 dmmu0.page_table\[5\]\[7\] net1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input252_I dcache_wb_adr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold288 dmmu1.page_table\[15\]\[1\] net1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold299 dmmu1.page_table\[12\]\[3\] net1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3936__S0 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3408_ _0875_ _1148_ _1149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7176_ net389 net642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4388_ _1956_ _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4884__I _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6127_ net200 _2974_ _2976_ dmmu1.page_table\[0\]\[12\] _2990_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3339_ _1069_ _1080_ _1081_ _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6058_ _2951_ _0516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5009_ _2265_ _2337_ _2339_ net759 _2341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6007__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2065 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4018__B1 _1669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4569__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_38_core_clock clknet_3_3_0_core_clock clknet_leaf_38_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5766__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5230__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3241__A1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_2082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5297__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7170__I net169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5049__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_77_core_clock clknet_3_5_0_core_clock clknet_leaf_77_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4257__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3359__B _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5509__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4980__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3690_ _1337_ net232 _1362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4732__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5360_ _2531_ _2535_ _2537_ net827 _2549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4311_ _1912_ _1910_ _1913_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5291_ _1808_ _2502_ _2504_ immu_0.page_table\[0\]\[5\] _2509_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_10_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7030_ net386 net408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4242_ net209 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3299__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4173_ _1812_ _1792_ _1794_ immu_0.page_table\[11\]\[6\] _1813_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7080__I net333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3124_ dmmu0.page_table\[8\]\[0\] dmmu0.page_table\[9\]\[0\] dmmu0.page_table\[10\]\[0\]
+ dmmu0.page_table\[11\]\[0\] _0872_ _0868_ _0874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_78_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3055_ net225 _0822_ _0828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_26_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1897 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6814_ _0387_ clknet_leaf_43_core_clock dmmu1.page_table\[11\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5748__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5212__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3223__A1 _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6745_ _0318_ clknet_leaf_39_core_clock dmmu1.page_table\[15\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3957_ _1618_ _1619_ _1416_ _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6676_ _0249_ clknet_leaf_34_core_clock dmmu0.page_table\[2\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3888_ net5 immu_0.high_addr_off\[0\] _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_33_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5627_ _2703_ _0333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6932__CLK clknet_leaf_58_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_2478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5558_ _2662_ _0305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_1201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input63_I c0_o_req_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4509_ _1909_ _2028_ _2031_ _2032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_28_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5489_ _2527_ _2613_ _2615_ dmmu0.page_table\[4\]\[8\] _2624_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_6_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4487__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7159_ net173 net629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_1565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6312__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5987__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3462__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6462__CLK clknet_leaf_99_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5203__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3907__B _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7165__I net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4714__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5911__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_1975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5690__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6805__CLK clknet_leaf_68_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__A2 _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4650__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4860_ _1797_ _2242_ _2244_ dmmu0.page_table\[9\]\[1\] _2246_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_1701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3811_ _1474_ immu_1.page_table\[15\]\[2\] _1479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6955__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4791_ _2203_ _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_17 net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6530_ _0103_ clknet_leaf_1_core_clock immu_0.page_table\[8\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3742_ immu_1.page_table\[8\]\[0\] immu_1.page_table\[9\]\[0\] immu_1.page_table\[10\]\[0\]
+ immu_1.page_table\[11\]\[0\] _1409_ _1410_ _1412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3300__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6155__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6461_ _0034_ clknet_leaf_11_core_clock dmmu0.page_table\[9\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7075__I net359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3673_ _1301_ _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_31_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5412_ immu_0.high_addr_off\[6\] _1812_ _2572_ _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6392_ _0774_ clknet_leaf_94_core_clock immu_1.page_table\[10\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5343_ _2540_ _0212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_71_2331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_46_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_2353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6335__CLK clknet_leaf_75_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5274_ _2498_ _0185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4469__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4225_ _1855_ _1841_ _1843_ immu_1.page_table\[9\]\[4\] _1856_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5130__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__I net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4156_ _1799_ _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3692__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6485__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3119__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3107_ net46 net45 net48 net47 _0857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_74_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_2271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5969__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_2282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4087_ net12 immu_0.high_addr_off\[7\] _1745_ _1746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_39_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input215_I dcache_mem_o_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_2293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3038_ _0812_ _0814_ _0816_ net603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_65_2146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5197__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4989_ _2327_ _0071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinterconnect_inner_712 c0_i_core_int_sreg[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_19_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinterconnect_inner_723 c1_i_core_int_sreg[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4944__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6728_ _0301_ clknet_leaf_41_core_clock dmmu0.page_table\[3\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4944__B2 dmmu0.page_table\[7\]\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_inner_734 c1_i_irq vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_22_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6659_ _0232_ clknet_leaf_23_core_clock dmmu0.page_table\[11\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_1105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput680 net680 inner_wb_adr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput691 net691 inner_wb_o_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output434_I net434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3358__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6828__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3181__C _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5672__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3683__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4880__B1 _2243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5424__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6978__CLK clknet_leaf_103_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3435__A1 _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3986__A2 _1647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6208__CLK clknet_leaf_73_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4935__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4935__B2 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput15 c0_o_mem_addr[11] net15 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 c0_o_mem_addr[7] net26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput37 c0_o_mem_data[2] net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput48 c0_o_mem_high_addr[3] net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput59 c0_o_req_addr[0] net59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6358__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5360__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3910__A2 _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5112__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4010_ _1670_ _1671_ _1367_ _1672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3674__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6175__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5961_ _2788_ _2890_ _2892_ dmmu1.page_table\[5\]\[4\] _2897_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4912_ _2278_ _0043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5892_ _2857_ _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_60_2010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4843_ _1817_ _2224_ _2226_ dmmu0.page_table\[10\]\[8\] _2235_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4774_ _1797_ _2191_ _2193_ immu_0.page_table\[12\]\[1\] _2195_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_56_894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6513_ _0086_ clknet_leaf_2_core_clock immu_0.page_table\[10\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3725_ _1370_ immu_0.page_table\[6\]\[0\] _1391_ _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6444_ _0017_ clknet_leaf_22_core_clock dmmu0.page_table\[10\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_2404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3656_ _1302_ net372 _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6375_ _0757_ clknet_leaf_78_core_clock immu_1.page_table\[11\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3587_ net215 _1219_ _1294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input165_I c1_o_req_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5326_ net104 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_3_2_0_core_clock clknet_0_core_clock clknet_3_2_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5103__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5257_ _1796_ _2486_ _2488_ immu_0.page_table\[1\]\[1\] _2490_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input332_I ic1_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4208_ _1842_ _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_3_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5188_ _1776_ _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3665__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input26_I c0_o_mem_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4862__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_2208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4892__I _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_2219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ net90 _1782_ _1784_ _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_19_1707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3760__S1 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3417__A1 net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_2034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4090__A1 net117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4917__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6500__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6119__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4132__I net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5342__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6650__CLK clknet_leaf_10_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5893__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3656__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3408__A1 _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4081__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4908__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5581__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3510_ net156 dmmu1.long_off_reg\[6\] _1248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4490_ _2020_ _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3441_ net49 dmmu0.long_off_reg\[4\] _1181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6160_ _3010_ _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3372_ _0938_ _1113_ _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5111_ _2399_ _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6091_ _2849_ _2958_ _2960_ net868 _2970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_40_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5097__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5636__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5042_ _2359_ _0092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3742__S1 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6993_ _0566_ clknet_leaf_94_core_clock dmmu1.long_off_reg\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_1339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6061__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3121__I _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5944_ _2886_ _0467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4072__A1 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_24_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6523__CLK clknet_leaf_2_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5875_ _2846_ _0438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_2051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4826_ _2225_ _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_12_2084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5021__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4375__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4757_ _1812_ _2175_ _2177_ net976 _2184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6673__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input282_I ic0_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3708_ _1377_ _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_43_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_1435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4688_ _2051_ _2139_ _2142_ net923 _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5324__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6427_ _0000_ clknet_leaf_105_core_clock immu_0.page_table\[13\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4127__A2 _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4887__I _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3639_ _0812_ net261 _1323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_1700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3335__B1 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6358_ _0740_ clknet_leaf_77_core_clock immu_1.page_table\[13\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3886__A1 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ _2451_ _2516_ _2518_ net820 _2520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput205 c1_sr_bus_data_o[5] net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6289_ _0671_ clknet_leaf_97_core_clock dmmu0.page_table\[0\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput216 dcache_mem_o_data[11] net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput227 dcache_mem_o_data[7] net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput238 dcache_wb_adr[16] net238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput249 dcache_wb_adr[4] net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4835__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4063__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5563__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5315__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7173__I net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5866__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3877__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5618__A2 _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3629__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold4 immu_0.page_table\[0\]\[0\] net738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_55_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6546__CLK clknet_leaf_3_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6043__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ net114 immu_1.high_addr_off\[4\] _1652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_69_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6696__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5660_ dmmu0.long_off_reg\[4\] _1806_ _2716_ _2721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ _2061_ _2090_ _2092_ immu_1.page_table\[13\]\[3\] _2096_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4357__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5591_ _1769_ _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_53_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4542_ _1838_ _1874_ _2028_ _2052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_68_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4109__A2 net255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ net208 _1999_ _2001_ immu_1.page_table\[1\]\[8\] _2010_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_20_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6212_ _0594_ clknet_leaf_94_core_clock immu_1.page_table\[9\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3424_ dmmu1.page_table\[0\]\[9\] dmmu1.page_table\[1\]\[9\] dmmu1.page_table\[2\]\[9\]
+ dmmu1.page_table\[3\]\[9\] _0886_ _0900_ _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3868__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3868__B2 net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6143_ _1980_ _2999_ _3001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3355_ _0938_ _1097_ _0879_ _1098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3116__I net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6074_ _2961_ _0522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3286_ dmmu0.page_table\[15\]\[4\] _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5025_ _2330_ _2337_ _2339_ immu_0.page_table\[10\]\[9\] _2349_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4293__A1 _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input128_I c1_o_mem_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_28_core_clock clknet_3_3_0_core_clock clknet_leaf_28_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_0_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__A1 net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6976_ _0549_ clknet_leaf_102_core_clock mem_dcache_arb.req1_pending vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__B2 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5242__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5927_ _2784_ _2873_ _2875_ net1057 _2878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5858_ _2682_ _2835_ _2837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_5_1281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input93_I c0_sr_bus_data_o[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _2215_ _0003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5545__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5789_ _2797_ _0401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6419__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5848__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3859__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Right_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_67_core_clock clknet_3_6_0_core_clock clknet_leaf_67_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4808__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output514_I net514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3706__S1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5481__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_1979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6025__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4036__A1 net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4587__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5784__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7168__I net167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4339__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_2077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3645__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_2039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput509 net509 c1_i_req_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_10_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4511__A2 _2032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Right_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3140_ net155 net154 net157 net156 _0890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_78_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3071_ _0836_ net470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4275__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4990__I net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6183__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _0403_ clknet_leaf_42_core_clock dmmu1.page_table\[10\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5775__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6761_ _0334_ clknet_leaf_31_core_clock dmmu0.page_table\[5\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3973_ _1631_ _1634_ _1635_ _1636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_53_Right_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7078__I net362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5712_ _2065_ _2743_ _2745_ net886 _2751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6692_ _0265_ clknet_leaf_91_core_clock immu_1.high_addr_off\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5527__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5643_ _2711_ _0341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5574_ _2672_ _0311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4525_ _1861_ _2033_ _2035_ dmmu1.page_table\[14\]\[6\] _2042_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold201 dmmu1.page_table\[2\]\[5\] net935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold212 immu_0.page_table\[14\]\[0\] net946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold223 dmmu1.page_table\[8\]\[0\] net957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5326__I net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold234 dmmu0.page_table\[2\]\[5\] net968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3274__C _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold245 dmmu0.page_table\[2\]\[12\] net979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ _2000_ _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xhold256 dmmu0.page_table\[8\]\[10\] net990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold267 immu_1.page_table\[11\]\[5\] net1001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_62_Right_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_103_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold278 immu_1.page_table\[8\]\[0\] net1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6711__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold289 dmmu0.page_table\[6\]\[7\] net1023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3407_ dmmu0.page_table\[4\]\[9\] dmmu0.page_table\[5\]\[9\] dmmu0.page_table\[6\]\[9\]
+ dmmu0.page_table\[7\]\[9\] _0871_ _0866_ _1148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7175_ net211 net639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3936__S1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4387_ _1839_ _1873_ _1909_ _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_input245_I dcache_wb_adr[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6126_ _2989_ _0546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3338_ net151 dmmu1.long_off_reg\[1\] _1081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6057_ _2794_ _2941_ _2943_ net918 _2951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3269_ net1 _1014_ _1015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6861__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5008_ _2340_ _0077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6007__A2 _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_71_Right_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5215__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_2090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5766__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4569__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ _0532_ clknet_leaf_62_core_clock dmmu1.page_table\[1\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_53_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3872__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6241__CLK clknet_leaf_93_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_80_Right_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4140__I net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6391__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output631_I net631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3552__I0 net138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4257__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5206__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_2076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5509__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4980__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3375__B _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6734__CLK clknet_leaf_44_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4732__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4310_ _1770_ _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_11_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5290_ _2508_ _0191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4241_ _1867_ _0592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_1179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3299__A2 _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6884__CLK clknet_leaf_48_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4040__S0 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_7_0_core_clock clknet_0_core_clock clknet_3_7_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4172_ _1811_ _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_78_1545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3123_ dmmu0.page_table\[12\]\[0\] dmmu0.page_table\[13\]\[0\] dmmu0.page_table\[14\]\[0\]
+ dmmu0.page_table\[15\]\[0\] _0872_ _0868_ _0873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_3054_ _0827_ net477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_1106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6813_ _0386_ clknet_leaf_41_core_clock dmmu1.page_table\[11\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5748__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6264__CLK clknet_leaf_84_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3956_ immu_1.page_table\[4\]\[7\] immu_1.page_table\[5\]\[7\] immu_1.page_table\[6\]\[7\]
+ immu_1.page_table\[7\]\[7\] _1404_ _1540_ _1619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6744_ _0317_ clknet_leaf_40_core_clock dmmu1.page_table\[15\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_63_2096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3223__A2 _0961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6675_ _0248_ clknet_leaf_33_core_clock dmmu0.page_table\[2\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3887_ _1422_ _1546_ _1551_ _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_45_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5626_ _1796_ _2699_ _2701_ dmmu0.page_table\[5\]\[1\] _2703_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input195_I c1_sr_bus_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5557_ net95 _2646_ _2648_ dmmu0.page_table\[3\]\[12\] _2662_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_2479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input362_I ic1_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4508_ _2030_ _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_13_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5488_ _2623_ _0274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input56_I c0_o_mem_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4895__I _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4439_ _1815_ _1979_ _1982_ dmmu0.page_table\[0\]\[7\] _1990_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4487__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5684__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7158_ net172 net628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6109_ _1851_ _2975_ _2977_ dmmu1.page_table\[0\]\[3\] _2981_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7089_ net343 net496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5436__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5987__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3837__I1 immu_1.page_table\[9\]\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6607__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3240__S _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1004 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4411__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6757__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output679_I net679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4962__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4714__A2 _2156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5911__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7181__I net400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3525__I0 net134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6287__CLK clknet_leaf_36_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4650__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3810_ _1405_ immu_1.page_table\[14\]\[2\] _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ _1819_ _2191_ _2193_ immu_0.page_table\[12\]\[9\] _2203_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_1735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_18 net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3741_ immu_1.page_table\[0\]\[0\] immu_1.page_table\[1\]\[0\] immu_1.page_table\[2\]\[0\]
+ immu_1.page_table\[3\]\[0\] _1409_ _1410_ _1411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_15_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6460_ _0033_ clknet_leaf_98_core_clock dmmu0.page_table\[9\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6155__A1 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3672_ _1345_ _1346_ _1347_ net680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_1470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5411_ _2578_ _0242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6391_ _0773_ clknet_leaf_77_core_clock immu_1.page_table\[10\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5342_ _2451_ _2536_ _2538_ dmmu0.page_table\[15\]\[1\] _2540_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_71_2332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5273_ net104 _2486_ _2488_ immu_0.page_table\[1\]\[9\] _2498_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4469__A1 _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4013__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4224_ _1854_ _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5130__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3141__A1 net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4155_ net97 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3692__A2 net365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3106_ net50 net49 net52 net51 _0856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_74_1217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _1744_ _1712_ _1745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5969__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_2272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6091__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3037_ net388 _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XTAP_TAPCELL_ROW_65_2147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input110_I c1_o_instr_long_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_2158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input208_I c1_sr_bus_data_o[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_2169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3995__S _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5197__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4988_ _2277_ _2317_ _2319_ net832 _2327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinterconnect_inner_713 c0_i_core_int_sreg[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_74_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_inner_724 c1_i_core_int_sreg[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_34_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6727_ _0300_ clknet_leaf_33_core_clock dmmu0.page_table\[3\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4944__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3939_ _1440_ _1602_ _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_22_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6658_ _0231_ clknet_leaf_28_core_clock dmmu0.page_table\[11\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_1909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4157__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5609_ _2692_ _0326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6589_ _0162_ clknet_leaf_17_core_clock immu_0.page_table\[3\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3235__S _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput670 net670 inner_wb_adr[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput681 net681 inner_wb_adr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput692 net692 inner_wb_o_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_79_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1964 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_1704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3034__I _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4880__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3683__A2 net378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4632__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4935__A2 _2290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7176__I net389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 c0_o_mem_addr[12] net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput27 c0_o_mem_addr[8] net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput38 c0_o_mem_data[3] net38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput49 c0_o_mem_high_addr[4] net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5360__A2 _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3653__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5112__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3674__A2 net376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6073__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5960_ _2896_ _0473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4911_ _2277_ _2261_ _2263_ net1056 _2278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5891_ _2682_ _2855_ _2857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_2000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_2022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4842_ _2234_ _0017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4926__A2 _2137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4773_ _2194_ _0797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6512_ _0085_ clknet_leaf_2_core_clock immu_0.page_table\[10\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3724_ _1385_ immu_0.page_table\[7\]\[0\] _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_67_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_2530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6302__CLK clknet_leaf_93_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3655_ _1332_ _1333_ _1334_ net676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6443_ _0016_ clknet_leaf_14_core_clock dmmu0.page_table\[10\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_2405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6374_ _0756_ clknet_leaf_72_core_clock immu_1.page_table\[11\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3586_ _1293_ net426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3362__A1 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5325_ _2528_ _0206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_1986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6452__CLK clknet_leaf_21_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input158_I c1_o_mem_long_mode vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5103__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5256_ _2489_ _0176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4207_ _1771_ _1840_ _1842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_3_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5187_ _2443_ _0153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3665__A2 net374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4862__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_2209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4138_ net82 net81 _1783_ _1784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_3_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input19_I c0_o_mem_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4069_ _1684_ _1727_ _1728_ _1729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4917__A2 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6119__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5342__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3353__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6945__CLK clknet_leaf_62_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3656__A2 net372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6055__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5802__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6325__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4908__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5419__I _2583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5581__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6475__CLK clknet_leaf_99_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3440_ net50 dmmu0.long_off_reg\[5\] _1180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3371_ dmmu0.page_table\[0\]\[8\] dmmu0.page_table\[1\]\[8\] dmmu0.page_table\[2\]\[8\]
+ dmmu0.page_table\[3\]\[8\] _0872_ _0941_ _1113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_21_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5110_ _2140_ _2397_ _2399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6090_ _2969_ _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_108_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5097__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5041_ _2271_ _2352_ _2354_ net1031 _2359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4993__I net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ _0565_ clknet_leaf_94_core_clock dmmu1.long_off_reg\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_18_core_clock clknet_3_2_0_core_clock clknet_leaf_18_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5943_ _2851_ _2872_ _2874_ net779 _2886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5874_ _2794_ _2836_ _2838_ net741 _2846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4825_ _1980_ _2223_ _2225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_47_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5021__A1 _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5329__I net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_58_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6818__CLK clknet_leaf_67_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4756_ _2183_ _0791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3583__A1 net228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4780__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3707_ net315 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4687_ _2141_ _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input275_I dcache_wb_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6426_ _0808_ clknet_leaf_106_core_clock immu_0.page_table\[13\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3638_ _1322_ net689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5324__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3335__A1 _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6968__CLK clknet_leaf_57_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3335__B2 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3569_ net221 _1204_ _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6357_ _0739_ clknet_leaf_76_core_clock immu_1.page_table\[13\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5308_ _2519_ _0198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6288_ _0670_ clknet_leaf_38_core_clock dmmu0.page_table\[0\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput206 c1_sr_bus_data_o[6] net206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_57_core_clock clknet_3_7_0_core_clock clknet_leaf_57_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput217 dcache_mem_o_data[12] net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput228 dcache_mem_o_data[8] net228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput239 dcache_wb_adr[17] net239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5239_ _2478_ _0170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4835__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_110_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output494_I net494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6498__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_49_Left_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5563__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output661_I net661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_96_core_clock clknet_3_4_0_core_clock clknet_leaf_96_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_34_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5315__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3326__A1 net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_60_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5079__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3629__A2 net271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold5 dmmu0.page_table\[12\]\[5\] net739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_37_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5251__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4610_ _2095_ _0733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5590_ _2680_ _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_26_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3565__A1 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4541_ _1823_ _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_20_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4472_ _2009_ _0681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3317__A1 net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6211_ _0593_ clknet_leaf_78_core_clock immu_1.page_table\[9\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3423_ _0896_ _1163_ _1164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7191_ net395 net648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3868__A2 _1532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6142_ _2999_ _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3354_ dmmu0.page_table\[0\]\[7\] dmmu0.page_table\[1\]\[7\] dmmu0.page_table\[2\]\[7\]
+ dmmu0.page_table\[3\]\[7\] _0950_ _0952_ _1097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6073_ _2776_ _2958_ _2960_ dmmu1.page_table\[1\]\[0\] _2961_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3285_ _0948_ _1027_ _1030_ _0940_ _1031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_77_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3176__S0 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5024_ _2348_ _0085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6019__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4293__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4228__I _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3132__I _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6975_ _0548_ clknet_leaf_102_core_clock mem_dcache_arb.select vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5242__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5926_ _2877_ _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6640__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5857_ _2835_ _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_75_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input392_I inner_wb_i_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _1806_ _2208_ _2210_ net831 _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5545__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5788_ _2103_ _2778_ _2780_ net782 _2797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input86_I c0_sr_bus_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4898__I _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6790__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4753__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4739_ _2171_ net76 _2172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_27_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6409_ _0791_ clknet_leaf_108_core_clock immu_0.page_table\[14\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3859__A2 _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5481__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_2025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output507_I net507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5784__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7184__I net403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6513__CLK clknet_leaf_2_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3070_ net217 _0831_ _0836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6663__CLK clknet_leaf_100_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5224__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6760_ _0333_ clknet_leaf_46_core_clock dmmu0.page_table\[5\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5775__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3972_ _1631_ _1634_ net2 _1635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3330__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5711_ _2750_ _0370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6691_ _0264_ clknet_leaf_89_core_clock immu_1.high_addr_off\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5642_ _2529_ _2699_ _2701_ dmmu0.page_table\[5\]\[9\] _2711_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5527__A2 _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3836__B _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ _2065_ _2664_ _2666_ dmmu1.page_table\[15\]\[5\] _2672_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4524_ _2041_ _0701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold202 dmmu1.page_table\[15\]\[9\] net936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_14_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold213 immu_0.page_table\[10\]\[2\] net947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold224 dmmu0.page_table\[3\]\[3\] net958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold235 dmmu0.page_table\[3\]\[6\] net969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold246 dmmu1.page_table\[11\]\[1\] net980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4455_ _1895_ _1998_ _2000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold257 immu_1.page_table\[4\]\[6\] net991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold268 dmmu1.page_table\[10\]\[7\] net1002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold279 dmmu1.page_table\[8\]\[6\] net1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6193__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3406_ _1145_ _1146_ _0877_ _1147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4386_ _1955_ _0649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7174_ net163 net638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3337_ net151 dmmu1.long_off_reg\[1\] _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6125_ net199 _2974_ _2976_ net1018 _2989_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_8_core_clock clknet_3_1_0_core_clock clknet_leaf_8_core_clock vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input140_I c1_o_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input238_I dcache_wb_adr[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3268_ net53 _1014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6056_ _2950_ _0515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5007_ _2258_ _2337_ _2339_ net899 _2340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3199_ _0867_ _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_55_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5215__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5766__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6958_ _0531_ clknet_leaf_62_core_clock dmmu1.page_table\[1\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_104_core_clock clknet_3_1_0_core_clock clknet_leaf_104_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_1377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3321__S0 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4974__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5909_ _2847_ _2856_ _2858_ dmmu1.page_table\[7\]\[8\] _2867_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6889_ _0462_ clknet_leaf_54_core_clock dmmu1.page_table\[6\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3872__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4726__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4421__I _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6536__CLK clknet_leaf_100_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output457_I net457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5453__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3388__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5151__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3552__I1 net33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6686__CLK clknet_leaf_92_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4257__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7179__I net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5206__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3768__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3312__S0 _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5509__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5390__B1 _2554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3940__A1 _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ _1866_ _1841_ _1843_ immu_1.page_table\[9\]\[8\] _1867_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4040__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4171_ net101 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3122_ _0871_ _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3053_ net224 _0822_ _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_26_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__CLK clknet_leaf_108_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6812_ _0385_ clknet_leaf_49_core_clock dmmu1.page_table\[11\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5748__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6743_ _0316_ clknet_leaf_39_core_clock dmmu1.page_table\[15\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4956__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_2086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3955_ immu_1.page_table\[0\]\[7\] immu_1.page_table\[1\]\[7\] immu_1.page_table\[2\]\[7\]
+ immu_1.page_table\[3\]\[7\] _1404_ _1540_ _1618_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_46_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_2097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6674_ _0247_ clknet_leaf_36_core_clock dmmu0.page_table\[2\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3886_ net107 _1549_ _1550_ _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6559__CLK clknet_leaf_4_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5625_ _2702_ _0332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5337__I _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input188_I c1_sr_bus_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3285__C _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5556_ _2661_ _0304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4507_ _1769_ _1837_ _2029_ _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_0_41_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5487_ _2463_ _2613_ _2615_ net1049 _2623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input355_I ic1_mem_data[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4438_ _1989_ _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4487__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5684__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I c0_o_mem_high_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7157_ net171 net627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4369_ _1849_ _1942_ _1944_ net776 _1947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6108_ _2980_ _0537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7088_ net341 net494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5436__A1 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6039_ _1891_ _1909_ _2030_ _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_9_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5987__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5372__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5911__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3922__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5124__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4650__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6701__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_19 net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3740_ net367 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_12_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6155__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3671_ _1337_ net251 _1347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5410_ immu_0.high_addr_off\[5\] _1809_ _2572_ _2578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6851__CLK clknet_leaf_36_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6390_ _0772_ clknet_leaf_80_core_clock immu_1.page_table\[10\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3913__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4996__I net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5341_ _2539_ _0211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_2333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5272_ _2497_ _0184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4013__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4469__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4223_ net204 _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3141__A2 net150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4154_ _1798_ _0574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5418__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3105_ _0855_ net519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6231__CLK clknet_leaf_83_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4085_ net11 immu_0.high_addr_off\[6\] _1744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5969__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_2273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6091__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_2284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3036_ _0812_ _0814_ _0815_ net602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_17_1603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_2148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4236__I _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input103_I c0_sr_bus_data_o[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6381__CLK clknet_leaf_72_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ _2326_ _0070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinterconnect_inner_714 c0_i_core_int_sreg[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_6726_ _0299_ clknet_leaf_35_core_clock dmmu0.page_table\[3\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3938_ immu_1.page_table\[0\]\[6\] immu_1.page_table\[1\]\[6\] immu_1.page_table\[2\]\[6\]
+ immu_1.page_table\[3\]\[6\] _1474_ _1433_ _1602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xinterconnect_inner_725 c1_i_core_int_sreg[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_22_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6657_ _0230_ clknet_leaf_14_core_clock dmmu0.page_table\[11\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3869_ inner_wb_arbiter.o_sel_sig _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_6_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4157__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5608_ _2463_ _2681_ _2684_ net1023 _2692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5354__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6588_ _0161_ clknet_leaf_14_core_clock immu_0.page_table\[3\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3904__A1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5539_ _2455_ _2647_ _2649_ net958 _2653_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput660 net660 inner_wb_adr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_2043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_54_1830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput671 net671 inner_wb_adr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput682 net682 inner_wb_adr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput693 net693 inner_wb_o_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_21_Left_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_35_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_65_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4880__A2 _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5530__I _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6724__CLK clknet_leaf_34_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3050__I _0825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Left_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6874__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput17 c0_o_mem_addr[13] net17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_1556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput28 c0_o_mem_addr[9] net28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput39 c0_o_mem_data[4] net39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5648__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6254__CLK clknet_leaf_84_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3754__S0 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_1505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5820__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4910_ _1814_ _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_73_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5890_ _2855_ _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_5_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_2001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _1815_ _2224_ _2226_ net1063 _2234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_60_2012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_2023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4387__A1 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4772_ _1777_ _2191_ _2193_ net1040 _2194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_16_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4926__A3 _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6511_ _0084_ clknet_leaf_0_core_clock immu_0.page_table\[10\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3723_ _1372_ _1388_ _1389_ _1392_ _1367_ _1393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_43_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_2520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_2531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6442_ _0015_ clknet_leaf_24_core_clock dmmu0.page_table\[10\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3654_ _1306_ net247 _1334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_73_2406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5887__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6373_ _0755_ clknet_leaf_72_core_clock immu_1.page_table\[11\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3585_ net229 _1219_ _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5324_ _2527_ _2516_ _2518_ net904 _2528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3993__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_47_core_clock clknet_3_6_0_core_clock clknet_leaf_47_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5255_ _1776_ _2486_ _2488_ immu_0.page_table\[1\]\[0\] _2489_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4311__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4206_ _1840_ _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_3_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5186_ _2332_ _2429_ _2431_ net878 _2443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4862__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4137_ net80 net79 net78 net77 _1783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA_input220_I dcache_mem_o_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input318_I ic0_wb_adr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4068_ net115 immu_1.high_addr_off\[5\] _1728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5662__I1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6897__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__I1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5575__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ _0282_ clknet_leaf_26_core_clock dmmu0.page_table\[13\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_1199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3976__I1 _1638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6119__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_86_core_clock clknet_3_5_0_core_clock clknet_leaf_86_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5327__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6277__CLK clknet_leaf_83_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput490 net490 c1_i_req_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5461__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6055__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5802__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7187__I net391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3041__A1 net559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3370_ _1110_ _1111_ _0938_ _1112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3975__S0 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5097__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5040_ _2358_ _0091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6991_ _0564_ clknet_leaf_94_core_clock dmmu1.long_off_reg\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5942_ _2885_ _0466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3280__A1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5873_ _2845_ _0437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4824_ _2223_ _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_7_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5021__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4755_ _1809_ _2175_ _2177_ immu_0.page_table\[14\]\[5\] _2183_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5309__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4780__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3583__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3706_ immu_0.page_table\[8\]\[0\] immu_0.page_table\[9\]\[0\] immu_0.page_table\[10\]\[0\]
+ immu_0.page_table\[11\]\[0\] _1370_ _1372_ _1376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_47_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4686_ _2140_ _2138_ _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6425_ _0807_ clknet_leaf_105_core_clock immu_0.page_table\[12\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3637_ _0812_ net260 _1322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_24_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input170_I c1_o_req_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input268_I dcache_wb_o_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3335__A2 _1076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6356_ _0738_ clknet_leaf_61_core_clock immu_1.page_table\[13\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3568_ _1284_ net411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5307_ _2444_ _2516_ _2518_ net1017 _2519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6287_ _0669_ clknet_leaf_36_core_clock dmmu0.page_table\[0\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3499_ dmmu0.page_table\[0\]\[12\] dmmu0.page_table\[1\]\[12\] dmmu0.page_table\[2\]\[12\]
+ dmmu0.page_table\[3\]\[12\] _0863_ _0866_ _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xinput207 c1_sr_bus_data_o[7] net207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput218 dcache_mem_o_data[13] net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput229 dcache_mem_o_data[9] net229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5238_ _2459_ _2470_ _2472_ net836 _2478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input31_I c0_o_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4835__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5169_ _2434_ _0144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6037__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4599__A1 _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output487_I net487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6912__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4523__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4523__B2 dmmu1.page_table\[14\]\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5720__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4287__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold6 immu_1.page_table\[8\]\[3\] net740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_76_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5539__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5003__A2 _2222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3565__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4540_ _2050_ _0708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6592__CLK clknet_leaf_4_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4471_ _1863_ _1999_ _2001_ immu_1.page_table\[1\]\[7\] _2009_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_1_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6210_ _0592_ clknet_leaf_79_core_clock immu_1.page_table\[9\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3422_ dmmu1.page_table\[4\]\[9\] dmmu1.page_table\[5\]\[9\] dmmu1.page_table\[6\]\[9\]
+ dmmu1.page_table\[7\]\[9\] _0886_ _0900_ _1163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7190_ net394 net647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6141_ _1826_ _1839_ _1892_ _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3353_ _0940_ _1095_ _1096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6072_ _2959_ _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3284_ _0882_ _1028_ _1029_ _0948_ _1030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_20_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5023_ _2328_ _2337_ _2339_ net992 _2348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3176__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6019__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5778__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6974_ _0547_ clknet_leaf_62_core_clock dmmu1.page_table\[0\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5242__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5925_ _2782_ _2873_ _2875_ net914 _2877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3253__A1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5856_ _1826_ _1892_ _2031_ _2835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XPHY_EDGE_ROW_3_Right_3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4807_ _2214_ _0002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5787_ _2796_ _0400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4753__A1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input385_I inner_embed_mode vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4738_ net83 _2171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_9_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input79_I c0_sr_bus_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4669_ _2130_ _0757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6408_ _0790_ clknet_leaf_107_core_clock immu_0.page_table\[14\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4505__A1 net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5702__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6339_ _0721_ clknet_leaf_75_core_clock immu_1.page_table\[14\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4269__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4808__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4419__I _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_2015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5481__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3492__A1 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5769__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4441__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3198__C _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5941__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_2079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6808__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_2017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3322__I2 dmmu1.page_table\[14\]\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3483__A1 _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6958__CLK clknet_leaf_62_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3971_ _1632_ _1633_ _1634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5710_ _2063_ _2743_ _2745_ dmmu1.page_table\[12\]\[4\] _2750_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6690_ _0263_ clknet_leaf_89_core_clock immu_1.high_addr_off\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3330__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1035 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5641_ _2710_ _0340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5572_ _2671_ _0310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4523_ _1858_ _2033_ _2035_ dmmu1.page_table\[14\]\[5\] _2041_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold203 immu_1.page_table\[6\]\[6\] net937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold214 dmmu1.page_table\[15\]\[4\] net948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_68_Left_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold225 dmmu1.page_table\[6\]\[8\] net959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4454_ _1998_ _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6338__CLK clknet_leaf_61_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold236 dmmu1.page_table\[4\]\[10\] net970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold247 dmmu1.page_table\[10\]\[0\] net981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4499__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold258 immu_0.page_table\[10\]\[8\] net992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold269 immu_0.page_table\[3\]\[2\] net1003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3405_ dmmu0.page_table\[8\]\[9\] dmmu0.page_table\[9\]\[9\] dmmu0.page_table\[10\]\[9\]
+ dmmu0.page_table\[11\]\[9\] _0871_ _0866_ _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_1_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7173_ net180 net637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4385_ _1870_ _1941_ _1943_ immu_1.page_table\[4\]\[10\] _1955_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3171__B1 _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6124_ _2988_ _0545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3336_ _1071_ _1079_ net526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__4239__I net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6488__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6055_ _2792_ _2941_ _2943_ net1059 _2950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3267_ net124 _0933_ _0989_ _1012_ _0841_ _1013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__5999__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input133_I c1_o_mem_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5006_ _2338_ _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_59_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3474__A1 _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3198_ _0879_ _0939_ _0946_ _0883_ _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XPHY_EDGE_ROW_77_Left_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input300_I ic0_mem_data[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5215__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_2081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6957_ _0530_ clknet_leaf_59_core_clock dmmu1.page_table\[1\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4974__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3321__S1 _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5908_ _2866_ _0451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6888_ _0461_ clknet_leaf_65_core_clock dmmu1.page_table\[6\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5839_ _2826_ _0422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4726__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5923__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5151__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3388__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3254__S _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4662__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5206__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3217__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3312__S1 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_72_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5390__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6630__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4170_ _1810_ _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3121_ _0863_ _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3052_ _0826_ net476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6780__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput390 inner_wb_i_dat[10] net390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_26_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6811_ _0384_ clknet_leaf_49_core_clock dmmu1.page_table\[11\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4405__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6742_ _0315_ clknet_leaf_66_core_clock dmmu1.page_table\[15\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4956__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3954_ net113 immu_1.high_addr_off\[3\] _1616_ _1617_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_63_2087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6673_ _0246_ clknet_leaf_37_core_clock dmmu0.page_table\[2\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3885_ _1547_ _1548_ _1550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5624_ _1776_ _2699_ _2701_ net797 _2702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4708__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5905__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5555_ net94 _2646_ _2648_ dmmu0.page_table\[3\]\[11\] _2661_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3138__I _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4506_ _1830_ net196 _1831_ _1832_ _2029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_13_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5486_ _2622_ _0273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4437_ _1812_ _1979_ _1982_ dmmu0.page_table\[0\]\[6\] _1989_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_6_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input250_I dcache_wb_adr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input348_I ic1_mem_data[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5684__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7156_ net164 net620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4368_ _1946_ _0640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6107_ _1848_ _2975_ _2977_ dmmu1.page_table\[0\]\[2\] _2980_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3319_ _1052_ _1063_ net525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7087_ net340 net493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4299_ _1863_ _1894_ _1897_ immu_1.page_table\[0\]\[7\] _1905_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_52_1780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5436__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6038_ _2939_ _0508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3447__A1 net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4644__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6503__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6149__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3249__S _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5372__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3048__I _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6653__CLK clknet_leaf_21_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5124__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3438__A1 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3670_ _0814_ net321 _1326_ _1346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5340_ _2444_ _2536_ _2538_ dmmu0.page_table\[15\]\[0\] _2539_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_51_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3913__A2 net239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5271_ net103 _2486_ _2488_ immu_0.page_table\[1\]\[8\] _2497_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xclkbuf_leaf_37_core_clock clknet_3_3_0_core_clock clknet_leaf_37_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_71_2334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4222_ _1853_ _0587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_1855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3677__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3141__A3 net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4153_ _1797_ _1792_ _1794_ immu_0.page_table\[11\]\[1\] _1798_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5418__A2 _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3104_ net119 net14 _0850_ _0855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4084_ _1306_ _1725_ _1742_ _1743_ net674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__3429__A1 _1154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_2274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6091__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_2285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3035_ net387 _0815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_37_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_2149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6526__CLK clknet_leaf_8_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4986_ _2275_ _2317_ _2319_ dmmu0.page_table\[14\]\[6\] _2326_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5051__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3937_ _1434_ _1600_ _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6725_ _0298_ clknet_leaf_13_core_clock dmmu0.page_table\[3\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinterconnect_inner_715 c0_i_core_int_sreg[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_inner_726 c1_i_core_int_sreg[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_73_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6676__CLK clknet_leaf_34_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input298_I ic0_mem_data[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6656_ _0229_ clknet_leaf_20_core_clock dmmu0.page_table\[11\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3868_ _1382_ _1532_ _1533_ net2 _1422_ _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xclkbuf_leaf_76_core_clock clknet_3_5_0_core_clock clknet_leaf_76_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_61_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5607_ _2691_ _0325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5354__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4157__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ _0160_ clknet_leaf_16_core_clock immu_0.page_table\[3\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3799_ _1375_ _1381_ _1466_ _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_15_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5538_ _2652_ _0295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input61_I c0_o_req_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_2011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5469_ _1976_ _2428_ _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_63_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput650 net650 ic1_wb_i_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput661 net661 inner_wb_adr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput672 net672 inner_wb_adr[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput683 net683 inner_wb_adr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput694 net694 inner_wb_o_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_50_1706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7139_ net211 net601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_6_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4617__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5459__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 c0_o_mem_addr[14] net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput29 c0_o_mem_data[0] net29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5648__A2 _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3203__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3659__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3754__S1 _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6549__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4084__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1946 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3831__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6699__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4840_ _2233_ _0016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_60_2002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3397__B _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _2192_ _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_16_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4387__A2 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6510_ _0083_ clknet_leaf_2_core_clock immu_0.page_table\[10\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3722_ _1385_ immu_0.page_table\[3\]\[0\] _1391_ _1392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_70_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_2510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6441_ _0014_ clknet_leaf_22_core_clock dmmu0.page_table\[10\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3653_ _0814_ net317 _1326_ _1333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_73_2407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6372_ _0754_ clknet_leaf_74_core_clock immu_1.page_table\[11\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3584_ _1292_ net425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_1944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3898__A1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5323_ net103 _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_12_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3993__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5254_ _2487_ _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4847__B1 _2225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4205_ _1829_ _1839_ _1840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5185_ _2442_ _0152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_3_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4136_ net91 _1782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_79_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4067_ net115 immu_1.high_addr_off\[5\] _1727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3151__I _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input213_I dcache_mem_exception vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_2037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5575__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4969_ _2315_ _0063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6708_ _0281_ clknet_leaf_25_core_clock dmmu0.page_table\[13\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5327__A1 _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6639_ _0212_ clknet_leaf_25_core_clock dmmu0.page_table\[15\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3527__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3889__A1 net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput480 net480 c1_i_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput491 net491 c1_i_req_data[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_output432_I net432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_1225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6055__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3061__I _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4066__A1 net116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6841__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5802__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3813__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5015__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_11_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6991__CLK clknet_leaf_94_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4106__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_2033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6221__CLK clknet_leaf_84_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3424__S0 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3975__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5652__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6371__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4829__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3680__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_2200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4057__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6990_ _0563_ clknet_leaf_102_core_clock inner_wb_arbiter.o_sel_sig vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__3104__I0 net119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5941_ _2849_ _2873_ _2875_ dmmu1.page_table\[6\]\[9\] _2885_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5872_ _2792_ _2836_ _2838_ net1013 _2845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _1977_ _2222_ _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_7_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5557__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4754_ _2182_ _0790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5309__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3705_ _1366_ _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4780__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4685_ _1770_ _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6424_ _0806_ clknet_leaf_107_core_clock immu_0.page_table\[12\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3636_ _1321_ net688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6714__CLK clknet_leaf_30_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6355_ _0737_ clknet_leaf_71_core_clock immu_1.page_table\[13\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3567_ net214 _1204_ _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3146__I net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1004 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input163_I c1_o_req_active vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5306_ _2517_ _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6286_ _0668_ clknet_leaf_33_core_clock dmmu0.page_table\[0\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3498_ net52 dmmu0.long_off_reg\[7\] _1235_ _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_52_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput208 c1_sr_bus_data_o[8] net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5237_ _2477_ _0169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput219 dcache_mem_o_data[14] net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_1460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6864__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input330_I ic1_mem_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_core_clock_I core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5168_ _2265_ _2430_ _2432_ net760 _2434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input24_I c0_o_mem_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6037__A2 _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4119_ _1772_ net462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4048__A1 net11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5099_ _2277_ _2382_ _2384_ immu_0.page_table\[7\]\[7\] _2392_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5796__A1 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_2_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6244__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_77_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3484__C _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6394__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4523__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5720__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4287__A1 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold7 dmmu1.page_table\[8\]\[7\] net741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_57_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4039__A1 net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5236__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3893__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5539__A1 _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6737__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4470_ _2008_ _0680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3421_ _1160_ _1161_ _0906_ _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6887__CLK clknet_leaf_52_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6140_ _2998_ _0551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3352_ dmmu0.page_table\[4\]\[7\] dmmu0.page_table\[5\]\[7\] dmmu0.page_table\[6\]\[7\]
+ dmmu0.page_table\[7\]\[7\] _0882_ _0948_ _1095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6071_ _1770_ _2957_ _2959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3283_ _0865_ dmmu0.page_table\[8\]\[4\] _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5475__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5022_ _2347_ _0084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6019__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5778__A1 _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6973_ _0546_ clknet_leaf_58_core_clock dmmu1.page_table\[0\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6267__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5924_ _2876_ _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5855_ _2834_ _0430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _1803_ _2208_ _2210_ immu_0.page_table\[13\]\[3\] _2214_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5786_ _2101_ _2778_ _2780_ net813 _2796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4737_ _2170_ _0785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4753__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input280_I ic0_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input378_I ic1_wb_adr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4668_ _2063_ _2123_ _2125_ immu_1.page_table\[11\]\[4\] _2130_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6407_ _0789_ clknet_leaf_105_core_clock immu_0.page_table\[14\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3619_ _1308_ net266 _1313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4505__A2 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5702__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4599_ _1870_ _2074_ _2076_ immu_1.page_table\[14\]\[10\] _2088_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4061__S0 _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6338_ _0720_ clknet_leaf_61_core_clock immu_1.page_table\[14\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6269_ _0651_ clknet_leaf_84_core_clock immu_1.page_table\[6\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4269__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3540__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5769__A1 _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4441__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output597_I net597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5467__S _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5941__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Right_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5209__B1 _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4680__A1 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3970_ net8 immu_0.high_addr_off\[3\] _1633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5640_ _2527_ _2699_ _2701_ dmmu0.page_table\[5\]\[8\] _2710_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_1446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_22_Right_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5571_ _2063_ _2664_ _2666_ net948 _2671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ _2040_ _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold204 immu_0.page_table\[11\]\[2\] net938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold215 immu_1.page_table\[2\]\[6\] net949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_48_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold226 dmmu1.page_table\[9\]\[1\] net960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4453_ _1828_ _1838_ _1891_ _1998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
Xhold237 immu_0.page_table\[8\]\[3\] net971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4499__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4043__S0 _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold248 dmmu1.page_table\[1\]\[4\] net982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_61_1722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3546__I0 net135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold259 immu_1.page_table\[8\]\[9\] net993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_40_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3404_ dmmu0.page_table\[12\]\[9\] dmmu0.page_table\[13\]\[9\] dmmu0.page_table\[14\]\[9\]
+ dmmu0.page_table\[15\]\[9\] _0871_ _0867_ _1145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7172_ net109 net636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4384_ _1954_ _0648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3171__A1 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6123_ _2851_ _2974_ _2976_ net1070 _2988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3335_ _0862_ _1076_ _1078_ _0860_ _0884_ _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6054_ _2949_ _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_31_Right_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5999__A1 _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3266_ _0915_ _0994_ _0999_ _1004_ _1011_ _1012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_5005_ _2140_ _2336_ _2338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3197_ _0943_ _0945_ _0879_ _0946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__3474__A2 _1212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input126_I c1_o_mem_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6902__CLK clknet_leaf_54_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_2069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6956_ _0529_ clknet_leaf_58_core_clock dmmu1.page_table\[1\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_1201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5907_ _2794_ _2856_ _2858_ net849 _2866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4974__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6887_ _0460_ clknet_leaf_52_core_clock dmmu1.page_table\[6\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5838_ _1805_ _2819_ _2821_ net1086 _2826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input91_I c0_sr_bus_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5923__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _2784_ _2778_ _2780_ net922 _2785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3785__I0 net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_12_Left_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_2075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5151__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_2086 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6432__CLK clknet_leaf_108_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output512_I net512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4662__A1 _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6582__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_2002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4414__A1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3217__A2 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6167__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_1610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5390__A2 _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27_core_clock clknet_3_2_0_core_clock clknet_leaf_27_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4025__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5678__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5660__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3120_ dmmu0.page_table\[0\]\[0\] dmmu0.page_table\[1\]\[0\] dmmu0.page_table\[2\]\[0\]
+ dmmu0.page_table\[3\]\[0\] _0865_ _0868_ _0870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6925__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3051_ net223 _0822_ _0826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_26_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput380 ic1_wb_sel[0] net380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_1813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput391 inner_wb_i_dat[11] net391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6810_ _0383_ clknet_leaf_49_core_clock dmmu1.page_table\[11\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4405__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5602__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_2108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6741_ _0314_ clknet_leaf_42_core_clock dmmu1.page_table\[15\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3953_ _1613_ _1615_ _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_42_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4956__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_2088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3884_ _1547_ _1548_ _1549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6672_ _0245_ clknet_leaf_33_core_clock dmmu0.page_table\[2\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6305__CLK clknet_leaf_93_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_66_core_clock clknet_3_6_0_core_clock clknet_leaf_66_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4169__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5905__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5623_ _2700_ _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_42_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5554_ _2660_ _0303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4505_ net190 net189 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_44_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5485_ _2461_ _2613_ _2615_ net905 _2622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6455__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4436_ _1988_ _0666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6181__I1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3144__A1 net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4341__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4367_ _1846_ _1942_ _1944_ net880 _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7155_ net395 net610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input243_I dcache_wb_adr[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6106_ _2979_ _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3318_ _0862_ _1061_ _1062_ _0860_ _0884_ _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7086_ net339 net492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4298_ _1904_ _0612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_52_1770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_2002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6037_ net200 _2923_ _2925_ net823 _2939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3249_ dmmu1.page_table\[2\]\[4\] dmmu1.page_table\[3\]\[4\] _0908_ _0995_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4644__A1 _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_2068 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6939_ _0512_ clknet_leaf_51_core_clock dmmu1.page_table\[2\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4713__I _2156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6149__A1 _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_16_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5372__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3383__A1 net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output462_I net462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5124__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3135__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6085__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5832__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6328__CLK clknet_leaf_62_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4399__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6478__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5899__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3374__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4571__B1 _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3175__S _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_2471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5270_ _2496_ _0183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_2324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4323__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4221_ _1852_ _1841_ _1843_ immu_1.page_table\[9\]\[3\] _1853_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3677__A2 net252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4152_ _1796_ _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3141__A4 net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3103_ _0854_ net541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4083_ _1535_ net245 _1743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3702__I _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_2264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3034_ _0813_ _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_69_2275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4985_ _2325_ _0069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5051__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6724_ _0297_ clknet_leaf_34_core_clock dmmu0.page_table\[3\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3936_ immu_1.page_table\[4\]\[6\] immu_1.page_table\[5\]\[6\] immu_1.page_table\[6\]\[6\]
+ immu_1.page_table\[7\]\[6\] _1474_ _1433_ _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_18_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinterconnect_inner_716 c0_i_core_int_sreg[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_18_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_7_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_inner_727 c1_i_core_int_sreg[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_50_1286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6655_ _0228_ clknet_leaf_27_core_clock dmmu0.page_table\[11\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3867_ net5 immu_0.high_addr_off\[0\] _1533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3149__I _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input193_I c1_sr_bus_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5606_ _2461_ _2681_ _2684_ net801 _2691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5354__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6586_ _0159_ clknet_leaf_21_core_clock immu_0.page_table\[3\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3798_ _1372_ _1461_ _1465_ _1377_ _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_15_965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3365__A1 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5537_ _2453_ _2647_ _2649_ net811 _2652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3085__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input360_I ic1_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput640 net640 ic1_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5468_ _2611_ _0266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input54_I c0_o_mem_req vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput651 net651 ic1_wb_i_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_54_1821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput662 net662 inner_wb_adr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput673 net673 inner_wb_adr[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4419_ _1976_ _1977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_61_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput684 net684 inner_wb_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput695 net695 inner_wb_o_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5399_ _2571_ _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_26_1491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7138_ net58 net600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7069_ net331 net484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4617__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5814__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_48_1647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3768__B net705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput19 c0_o_mem_addr[15] net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_1812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6770__CLK clknet_leaf_38_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3203__S1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3659__A2 net248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4856__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_84_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4084__A2 _1725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_2003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5033__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_2014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _2140_ _2190_ _2192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4387__A3 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3595__A1 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3721_ _1390_ _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_15_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_2511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6440_ _0013_ clknet_leaf_28_core_clock dmmu0.page_table\[10\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_2533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3652_ _1302_ net371 _1332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_2012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3347__A1 _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_2408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3583_ net228 _1219_ _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6371_ _0753_ clknet_leaf_78_core_clock immu_1.page_table\[11\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5322_ _2526_ _0205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5253_ _1895_ _2485_ _2487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4847__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4204_ _1838_ _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5184_ _2330_ _2430_ _2432_ net1079 _2442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6049__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4135_ _1779_ _1780_ _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_3_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4066_ net116 immu_1.high_addr_off\[6\] _1726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_78_1197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6643__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input206_I c1_sr_bus_data_o[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4968_ _1996_ _2298_ _2301_ dmmu0.page_table\[7\]\[12\] _2315_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5575__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6707_ _0280_ clknet_leaf_25_core_clock dmmu0.page_table\[13\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3130__S0 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6793__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3919_ immu_0.page_table\[4\]\[6\] immu_0.page_table\[5\]\[6\] immu_0.page_table\[6\]\[6\]
+ immu_0.page_table\[7\]\[6\] _1424_ _1455_ _1583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_4899_ _2269_ _2261_ _2263_ net822 _2270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6638_ _0211_ clknet_leaf_25_core_clock dmmu0.page_table\[15\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5327__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3338__A1 net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6569_ _0142_ clknet_leaf_6_core_clock immu_0.page_table\[5\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput470 net470 c1_i_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput481 net481 c1_i_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput492 net492 c1_i_req_data[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3510__A1 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5263__A1 _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5015__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Right_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_26_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3577__A1 net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4901__I _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3424__S1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6516__CLK clknet_leaf_7_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_78_Right_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4829__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Left_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3188__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6666__CLK clknet_leaf_104_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_2201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3104__I1 net14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5940_ _2884_ _0465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5871_ _2844_ _0436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4822_ _1779_ _2172_ _2222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_70_1971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5557__A2 _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4016__C _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4753_ _1806_ _2175_ _2177_ net846 _2182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3704_ _1368_ _1373_ _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5309__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4684_ _2138_ _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_71_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6423_ _0805_ clknet_leaf_106_core_clock immu_0.page_table\[12\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4517__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3635_ _0812_ net259 _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6196__CLK clknet_leaf_108_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6354_ _0736_ clknet_leaf_75_core_clock immu_1.page_table\[13\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3566_ _1283_ net410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5305_ _2300_ _2515_ _2517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3497_ _1229_ _1233_ _1234_ _1235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6285_ _0667_ clknet_leaf_36_core_clock dmmu0.page_table\[0\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input156_I c1_o_mem_high_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput209 c1_sr_bus_data_o[9] net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5236_ _2457_ _2470_ _2472_ net1088 _2477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5493__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5167_ _2433_ _0143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3162__I net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input323_I ic0_wb_adr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4118_ icore_sregs.c1_disable net384 _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5098_ _2391_ _0116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input17_I c0_o_mem_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4049_ net10 immu_0.high_addr_off\[5\] _1709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_36_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5796__A2 _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3538__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6539__CLK clknet_leaf_3_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output542_I net542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4287__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4168__I _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold8 dmmu0.page_table\[5\]\[10\] net742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5236__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3098__I0 net131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_2044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3798__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3342__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4117__B _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3893__S1 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5539__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_971 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4747__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3970__A1 net8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ dmmu1.page_table\[8\]\[9\] dmmu1.page_table\[9\]\[9\] dmmu1.page_table\[10\]\[9\]
+ dmmu1.page_table\[11\]\[9\] _0887_ _0900_ _1161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5172__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_2037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1915 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_957 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3722__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3351_ net106 net158 _0884_ _1093_ _1094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_0_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6070_ _2957_ _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3282_ dmmu0.page_table\[9\]\[4\] _1028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5475__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I c0_o_instr_long_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5021_ _2277_ _2337_ _2339_ net891 _2347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3089__I0 net127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6972_ _0545_ clknet_leaf_62_core_clock dmmu1.page_table\[0\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5778__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5923_ _2776_ _2873_ _2875_ net756 _2876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4986__B1 _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5854_ net95 _2818_ _2820_ dmmu0.page_table\[1\]\[12\] _2834_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _2213_ _0001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5785_ _2795_ _0399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4541__I _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4736_ _1821_ _2156_ _2158_ net1027 _2170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3961__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4667_ _2129_ _0756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3157__I _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input273_I dcache_wb_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6406_ _0788_ clknet_leaf_110_core_clock immu_0.page_table\[14\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__CLK clknet_leaf_68_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3618_ _1312_ net694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5702__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ _2087_ _0729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4061__S1 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6337_ _0719_ clknet_leaf_71_core_clock immu_1.page_table\[15\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3549_ _1274_ net545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3093__S _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6268_ _0650_ clknet_leaf_82_core_clock immu_1.page_table\[6\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4269__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6981__CLK clknet_leaf_73_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5219_ _2330_ _2447_ _2449_ net870 _2466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6199_ _0581_ clknet_leaf_2_core_clock immu_0.page_table\[11\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6211__CLK clknet_leaf_78_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5769__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3324__S0 _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4441__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6361__CLK clknet_leaf_61_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output492_I net492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4044__I2 _1703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5941__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_core_clock clknet_3_2_0_core_clock clknet_leaf_17_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3704__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1093 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_23_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5209__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3530__I _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6704__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5658__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_56_core_clock clknet_3_7_0_core_clock clknet_leaf_56_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_80_2595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6854__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5570_ _2670_ _0309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4521_ _1855_ _2033_ _2035_ dmmu1.page_table\[14\]\[4\] _2040_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold205 immu_0.page_table\[3\]\[3\] net939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_79_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5145__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4452_ _1997_ _0673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold216 dmmu1.page_table\[1\]\[5\] net950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold227 immu_0.page_table\[9\]\[2\] net961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_48_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold238 immu_0.page_table\[9\]\[1\] net972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_65_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4499__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold249 immu_1.page_table\[7\]\[2\] net983 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_22_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4043__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5696__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3546__I1 net30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3403_ _1119_ _1143_ _1144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7171_ net170 net626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4383_ _1868_ _1942_ _1944_ immu_1.page_table\[4\]\[9\] _1954_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3705__I _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3171__A2 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6122_ _2987_ _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3334_ net46 dmmu0.long_off_reg\[1\] _1077_ _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_0_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5448__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6234__CLK clknet_leaf_93_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6053_ _2790_ _2941_ _2943_ net935 _2949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5920__I _2872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3265_ _0907_ _1007_ _1010_ _0912_ _1011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__5999__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4120__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5004_ _2336_ _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3196_ _0938_ _0944_ _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_95_core_clock clknet_3_4_0_core_clock clknet_leaf_95_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_18_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6384__CLK clknet_leaf_72_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input119_I c1_o_mem_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6955_ _0528_ clknet_leaf_56_core_clock dmmu1.page_table\[1\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5620__A1 _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4423__A2 _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5906_ _2865_ _0450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_1369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6886_ _0459_ clknet_leaf_49_core_clock dmmu1.page_table\[6\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5837_ _2825_ _0421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5367__I _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input390_I inner_wb_i_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5384__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5768_ _1848_ _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input84_I c0_sr_bus_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3934__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4719_ _2161_ _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5699_ _2742_ _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_20_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6727__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output505_I net505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_89_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4414__A2 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6877__CLK clknet_leaf_54_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6167__A2 net255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5277__I _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3925__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_955 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4025__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4102__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3050_ _0825_ net475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput370 ic1_wb_adr[1] net370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput381 ic1_wb_sel[1] net381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_26_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5850__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput392 inner_wb_i_dat[12] net392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_76_1284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5602__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4405__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5453__I1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6740_ _0313_ clknet_leaf_41_core_clock dmmu1.page_table\[15\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3952_ _1606_ _1549_ _1614_ _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_1408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6671_ _0244_ clknet_leaf_101_core_clock immu_0.high_addr_off\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3883_ net111 immu_1.high_addr_off\[1\] _1548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_50_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4169__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5622_ _2682_ _2698_ _2700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3216__I0 _0962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5905__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_868 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3916__A1 net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5553_ _2531_ _2646_ _2648_ dmmu0.page_table\[3\]\[10\] _2660_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_1954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_91_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4504_ _2027_ _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5118__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5484_ _2621_ _0272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4435_ _1809_ _1979_ _1982_ net884 _1988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_841 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4341__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7154_ net394 net609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4366_ _1945_ _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6105_ _1845_ _2975_ _2977_ dmmu1.page_table\[0\]\[1\] _2979_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3317_ net45 dmmu0.long_off_reg\[0\] _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7085_ net338 net491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4297_ _1860_ _1894_ _1897_ immu_1.page_table\[0\]\[6\] _1904_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_52_1760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input236_I dcache_wb_adr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _2938_ _0507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3248_ _0931_ _0990_ _0993_ _0906_ _0994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_33_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4644__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3179_ _0907_ _0927_ _0928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input403_I inner_wb_i_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6938_ _0511_ clknet_leaf_50_core_clock dmmu1.page_table\[2\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6149__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6869_ _0442_ clknet_leaf_66_core_clock dmmu1.page_table\[8\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_46_1597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3546__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3135__A2 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output622_I net622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5560__I _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3281__S _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6085__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3518__S0 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4176__I _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3080__I _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4904__I _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4399__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5596__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_7_core_clock clknet_3_0_0_core_clock clknet_leaf_7_core_clock vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_1165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5899__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4571__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_2450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4220_ _1851_ _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4323__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_103_core_clock clknet_3_1_0_core_clock clknet_leaf_103_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4874__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4151_ net96 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5470__I _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3102_ net133 net28 _0850_ _0854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4082_ _1422_ _1732_ _1741_ _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_21_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_69_2265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3033_ icache_arbiter.o_sel_sig _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_69_2276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ _2273_ _2317_ _2319_ dmmu0.page_table\[14\]\[5\] _2325_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5051__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_2097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6723_ _0296_ clknet_leaf_45_core_clock dmmu0.page_table\[3\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3062__A1 net228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3935_ _1502_ _1596_ _1598_ _1599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xinterconnect_inner_706 c0_i_core_int_sreg[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_34_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6422__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_inner_717 c0_i_core_int_sreg[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_inner_728 c1_i_core_int_sreg[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_74_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6654_ _0227_ clknet_leaf_27_core_clock dmmu0.page_table\[11\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3866_ _1525_ _1527_ _1529_ _1531_ _1532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_6_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5605_ _2690_ _0324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_41_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6585_ _0158_ clknet_leaf_16_core_clock immu_0.page_table\[3\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3797_ _1391_ _1462_ _1464_ _1465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_14_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input186_I c1_sr_bus_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3996__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5536_ _2651_ _0294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_1735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6572__CLK clknet_leaf_3_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5467_ immu_1.high_addr_off\[7\] _1864_ _2603_ _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3165__I net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput630 net630 ic1_mem_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput641 net641 ic1_wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input353_I ic1_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput652 net652 ic1_wb_i_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5511__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4418_ _1769_ _1788_ _1975_ _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_4
Xoutput663 net663 inner_wb_adr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput674 net674 inner_wb_adr[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5398_ _1785_ _2570_ _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input47_I c0_o_mem_high_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput685 net685 inner_wb_o_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput696 net696 inner_wb_o_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7137_ net75 net599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ _1858_ _1927_ _1929_ net1071 _1935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_35_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6067__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7068_ net407 net465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4617__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5814__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6019_ _2786_ _2924_ _2926_ net768 _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3053__A1 net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_1895 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3784__B _1452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6915__CLK clknet_leaf_54_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3276__S _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5750__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4305__A1 net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4856__A2 _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1890 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_2080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5656__I1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3816__B1 _1473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3292__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5408__I1 _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6445__CLK clknet_leaf_23_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5569__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_2004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5033__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_2015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5666__S _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3720_ net313 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_2095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3595__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4792__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6595__CLK clknet_leaf_21_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_2512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3651_ _1329_ _1330_ _1331_ net671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4544__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _0752_ clknet_leaf_70_core_clock immu_1.page_table\[12\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_2409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3582_ _1291_ net424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5321_ _2463_ _2516_ _2518_ net1084 _2526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ _2485_ _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4847__A2 _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4203_ _1769_ _1834_ _1837_ _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_4
XANTENNA__3713__I _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5183_ _2441_ _0151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6049__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4134_ net83 net76 _1780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_58_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1990 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4065_ _1712_ _1713_ _1718_ _1724_ _0813_ _1725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_56_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3283__A1 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input101_I c0_sr_bus_data_o[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6938__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4967_ _2314_ _0062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_43_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3130__S1 _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3918_ net7 immu_0.high_addr_off\[2\] _1581_ _1582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_30_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6706_ _0279_ clknet_leaf_69_core_clock dmmu0.page_table\[4\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4898_ _1802_ _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_69_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6637_ _0210_ clknet_leaf_10_core_clock dmmu0.page_table\[12\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3849_ immu_1.page_table\[12\]\[4\] immu_1.page_table\[13\]\[4\] immu_1.page_table\[14\]\[4\]
+ immu_1.page_table\[15\]\[4\] _1441_ _1442_ _1515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3096__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5732__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6568_ _0141_ clknet_leaf_4_core_clock immu_0.page_table\[5\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5519_ _2527_ _2630_ _2632_ net1024 _2641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_37_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6499_ _0072_ clknet_leaf_21_core_clock dmmu0.page_table\[14\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_37_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4299__B1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput460 net460 c0_i_req_data_valid vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput471 net471 c1_i_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput482 net482 c1_i_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput493 net493 c1_i_req_data[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_57_1205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_28_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3274__A1 _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5015__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1968 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4774__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3577__A2 _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5971__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1919 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4829__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3188__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_2202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3689__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3265__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5870_ _2790_ _2836_ _2838_ net847 _2844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4821_ _2221_ _0009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4752_ _2181_ _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4765__A1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3703_ immu_0.page_table\[12\]\[0\] immu_0.page_table\[13\]\[0\] immu_0.page_table\[14\]\[0\]
+ immu_0.page_table\[15\]\[0\] _1370_ _1372_ _1373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA_clkbuf_leaf_30_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4683_ _1839_ _2137_ _2138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3708__I _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6422_ _0804_ clknet_leaf_106_core_clock immu_0.page_table\[12\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4517__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3634_ _1320_ net687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4517__B2 dmmu1.page_table\[14\]\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5714__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5190__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6353_ _0735_ clknet_leaf_61_core_clock immu_1.page_table\[13\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3565_ net212 _1204_ _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_1874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5304_ _2515_ _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_59_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6284_ _0666_ clknet_leaf_38_core_clock dmmu0.page_table\[0\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3496_ net51 dmmu0.long_off_reg\[6\] _1234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_1077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5235_ _2476_ _0168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6610__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5493__A2 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input149_I c1_o_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5166_ _2258_ _2430_ _2432_ net882 _2433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4117_ _1764_ _1768_ _1771_ net684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_1536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ _2275_ _2382_ _2384_ immu_0.page_table\[7\]\[6\] _2391_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input316_I ic0_wb_adr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4048_ net11 immu_0.high_addr_off\[6\] _1708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3256__A1 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1080 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5999_ _2847_ _2907_ _2909_ dmmu1.page_table\[4\]\[8\] _2918_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_1411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5953__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3554__S _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3781__C _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6290__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3495__A1 net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4692__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold9 immu_0.page_table\[4\]\[8\] net743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_57_1013 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5236__A2 _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3247__A1 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3098__I1 net26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3342__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_46_core_clock clknet_3_6_0_core_clock clknet_leaf_46_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_1765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3528__I _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_2076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3972__B net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5172__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6633__CLK clknet_leaf_23_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_96_core_clock_I clknet_3_4_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_3350_ _0894_ _1083_ _1092_ _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3281_ dmmu0.page_table\[10\]\[4\] dmmu0.page_table\[11\]\[4\] _0865_ _1027_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5475__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5020_ _2346_ _0083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_85_core_clock clknet_3_5_0_core_clock clknet_leaf_85_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3089__I1 net22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4435__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6971_ _0544_ clknet_leaf_60_core_clock dmmu1.page_table\[0\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_928 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ _2874_ _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4986__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5853_ _2833_ _0429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4804_ _1800_ _2208_ _2210_ immu_0.page_table\[13\]\[2\] _2213_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5935__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5784_ _2794_ _2778_ _2780_ net1002 _2795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4202__A3 _1836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4735_ _2169_ _0784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3410__A1 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ _2061_ _2123_ _2125_ net844 _2129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6405_ _0787_ clknet_leaf_110_core_clock immu_0.page_table\[14\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3617_ _1308_ net265 _1312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4597_ _1868_ _2075_ _2077_ immu_1.page_table\[14\]\[9\] _2087_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input266_I dcache_wb_o_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6336_ _0718_ clknet_leaf_77_core_clock immu_1.page_table\[15\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3548_ net136 net31 _1267_ _1274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6267_ _0649_ clknet_leaf_87_core_clock immu_1.page_table\[4\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3479_ _1209_ _1214_ _1217_ _1051_ _1218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5218_ _2465_ _0162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6198_ _0580_ clknet_leaf_0_core_clock immu_0.page_table\[11\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4674__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5149_ _2273_ _2414_ _2416_ immu_0.page_table\[5\]\[5\] _2422_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3324__S1 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6506__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1096 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4044__I3 _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output485_I net485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6656__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4179__I net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6103__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4907__I _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_2009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5209__A2 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4968__A1 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_28_Left_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4520_ _2039_ _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold206 immu_1.page_table\[8\]\[6\] net940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4451_ _1996_ _1978_ _1981_ dmmu0.page_table\[0\]\[12\] _1997_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_1568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5145__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold217 immu_0.page_table\[5\]\[2\] net951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold228 immu_1.page_table\[10\]\[3\] net962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_65_1860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3402_ net49 dmmu0.long_off_reg\[4\] _1142_ _1143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5696__A2 _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold239 dmmu0.page_table\[15\]\[9\] net973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7170_ net169 net625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4382_ _1953_ _0647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3207__B _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6121_ _2849_ _2975_ _2977_ net966 _2987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_61_1757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3333_ net45 dmmu0.long_off_reg\[0\] _1077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_37_Left_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6052_ _2948_ _0513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_7_Right_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3459__A1 _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3264_ _0889_ _1008_ _1009_ _0931_ _1010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_77_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5003_ _1790_ _2222_ _2336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4120__A2 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3721__I _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3195_ dmmu0.page_table\[0\]\[1\] dmmu0.page_table\[1\]\[1\] dmmu0.page_table\[2\]\[1\]
+ dmmu0.page_table\[3\]\[1\] _0864_ _0867_ _0944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_20_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6529__CLK clknet_leaf_8_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6954_ _0527_ clknet_leaf_55_core_clock dmmu1.page_table\[1\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5905_ _2792_ _2856_ _2858_ dmmu1.page_table\[7\]\[6\] _2865_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3631__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ _0458_ clknet_leaf_52_core_clock dmmu1.page_table\[6\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6679__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_46_Left_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5836_ _1802_ _2819_ _2821_ dmmu0.page_table\[1\]\[3\] _2825_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5384__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5767_ _2783_ _0393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1960 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input383_I ic1_wb_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4718_ _1797_ _2157_ _2159_ immu_0.page_table\[15\]\[1\] _2161_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5698_ _1892_ _2028_ _2031_ _2742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_47_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input77_I c0_sr_bus_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4649_ _2118_ _0749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_1067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Left_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6319_ _0701_ clknet_leaf_96_core_clock dmmu1.page_table\[14\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4111__A2 net379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7103__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3870__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Left_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_1860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_1937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_923 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_1281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3481__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3806__I _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_73_Left_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_1129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5678__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3233__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3689__A1 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4102__A2 net326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3541__I _1270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput360 ic1_mem_data[7] net360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput371 ic1_wb_adr[2] net371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput382 ic1_wb_stb net382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5850__A2 _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput393 inner_wb_i_dat[13] net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3861__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6821__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5063__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5602__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3951_ net112 immu_1.high_addr_off\[2\] _1614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3613__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4810__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6670_ _0243_ clknet_leaf_101_core_clock immu_0.high_addr_off\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3882_ net110 immu_1.high_addr_off\[0\] _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5621_ _2698_ _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_73_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4169__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5552_ _2659_ _0302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4503_ _1870_ _2013_ _2015_ immu_1.page_table\[3\]\[10\] _2027_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5118__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5483_ _2459_ _2613_ _2615_ net799 _2621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6201__CLK clknet_leaf_100_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4434_ _1987_ _0665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3224__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7153_ net393 net608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4365_ _1824_ _1942_ _1944_ immu_1.page_table\[4\]\[0\] _1945_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4341__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6104_ _2978_ _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3316_ _1054_ _1056_ _1058_ _1060_ _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__6351__CLK clknet_leaf_75_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7084_ net337 net490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4296_ _1903_ _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_52_1761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6035_ net199 _2923_ _2925_ dmmu1.page_table\[3\]\[11\] _2938_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_52_1772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3247_ _0889_ _0991_ _0992_ _0902_ _0993_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_52_1783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input131_I c1_o_mem_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input229_I dcache_mem_o_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3178_ dmmu1.page_table\[0\]\[1\] dmmu1.page_table\[1\]\[1\] dmmu1.page_table\[2\]\[1\]
+ dmmu1.page_table\[3\]\[1\] _0888_ _0910_ _0927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_59_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6937_ _0510_ clknet_leaf_56_core_clock dmmu1.page_table\[2\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4282__I _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6868_ _0441_ clknet_leaf_66_core_clock dmmu1.page_table\[8\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_46_1587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_2081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5819_ _2814_ _0414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6799_ _0372_ clknet_leaf_50_core_clock dmmu1.page_table\[12\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3215__S0 _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4868__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output448_I net448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_1826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6085__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3518__S1 net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4096__A1 _1747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__CLK clknet_leaf_67_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5293__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5832__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3843__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5045__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5596__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4399__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6994__CLK clknet_leaf_95_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5899__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4020__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3454__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_35_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4571__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_2451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6374__CLK clknet_leaf_72_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_2326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4323__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_2348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ _1795_ _0573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3101_ _0853_ net540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4081_ _1502_ _1735_ _1740_ _1408_ _1741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4087__A1 net12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_2100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3032_ inner_wb_arbiter.o_sel_sig _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_69_2266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput190 c1_sr_bus_addr[3] net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_69_2277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1082 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4983_ _2324_ _0068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6722_ _0295_ clknet_leaf_36_core_clock dmmu0.page_table\[3\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3934_ _1434_ _1597_ _1598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3062__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_inner_707 c0_i_core_int_sreg[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_inner_718 c0_i_core_int_sreg[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_18_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinterconnect_inner_729 c1_i_core_int_sreg[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_15_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3865_ _1375_ _1530_ _1383_ _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6653_ _0226_ clknet_leaf_21_core_clock dmmu0.page_table\[11\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5604_ _2459_ _2681_ _2684_ dmmu0.page_table\[6\]\[5\] _2690_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_41_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3796_ _1463_ immu_0.page_table\[15\]\[2\] _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6584_ _0157_ clknet_leaf_14_core_clock immu_0.page_table\[3\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_1097 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6717__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5535_ _2451_ _2647_ _2649_ dmmu0.page_table\[3\]\[1\] _2651_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3996__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5466_ _2610_ _0265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input179_I c1_o_req_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput620 net620 ic1_mem_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_28_1769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput631 net631 ic1_mem_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput642 net642 ic1_wb_i_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4417_ _1974_ net91 _1784_ _1975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5511__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput653 net653 ic1_wb_i_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput664 net664 inner_wb_adr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5397_ _1895_ net105 _2569_ _2570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput675 net675 inner_wb_adr[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6867__CLK clknet_leaf_65_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput686 net686 inner_wb_o_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input346_I ic1_mem_data[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput697 net697 inner_wb_o_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4348_ _1934_ _0632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7136_ net4 net598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4277__I _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6067__A2 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7067_ net407 net464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4279_ net188 net181 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XANTENNA__5814__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6018_ _2929_ _0498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_1832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6247__CLK clknet_leaf_84_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3053__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6397__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3436__S0 _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output565_I net565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5750__A1 _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_2043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3816__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_2130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5569__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_2005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_2016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3650_ _1306_ net242 _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_77_2513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3581_ net227 _1204_ _1291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5320_ _2525_ _0204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_1936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5251_ _1789_ _2484_ _2485_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_45_1368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4202_ net210 _1835_ _1836_ _1837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5182_ _2328_ _2430_ _2432_ net743 _2441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6049__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4133_ _1778_ net84 _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_48_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5257__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4064_ _1382_ _1723_ _1724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5009__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_1115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4966_ _1994_ _2298_ _2301_ dmmu0.page_table\[7\]\[11\] _2314_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_43_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6705_ _0278_ clknet_leaf_38_core_clock dmmu0.page_table\[4\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3917_ _1553_ _1554_ _1580_ _1581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_46_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4897_ _2268_ _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4560__I _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input296_I ic0_mem_data[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6636_ _0209_ clknet_leaf_12_core_clock dmmu0.page_table\[12\]\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3848_ _1514_ net666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5732__A1 _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3779_ immu_1.page_table\[12\]\[1\] immu_1.page_table\[13\]\[1\] immu_1.page_table\[14\]\[1\]
+ immu_1.page_table\[15\]\[1\] _1441_ _1442_ _1448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_6567_ _0140_ clknet_leaf_18_core_clock immu_0.page_table\[5\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5518_ _2640_ _0287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6498_ _0071_ clknet_leaf_26_core_clock dmmu0.page_table\[14\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput450 net450 c0_i_req_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5449_ net191 _1836_ _2600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4299__A1 _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput461 net461 c0_rst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput472 net472 c1_i_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput483 net483 c1_i_mem_exception vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput494 net494 c1_i_req_data[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_61_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7119_ net395 net572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_3_5_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7111__I net402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4471__A1 _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36_core_clock clknet_3_3_0_core_clock clknet_leaf_36_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_26_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5420__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output682_I net682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4774__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5971__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3409__S0 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3086__I _0845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5487__B1 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6412__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3352__I3 dmmu0.page_table\[7\]\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_75_core_clock clknet_3_5_0_core_clock clknet_leaf_75_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_66_2203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6562__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4820_ _1821_ _2207_ _2209_ immu_0.page_table\[13\]\[10\] _2221_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_2084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4765__A2 _2174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4751_ _1803_ _2175_ _2177_ net1090 _2181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3702_ _1371_ _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4682_ _1826_ _1909_ _2137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_71_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6421_ _0803_ clknet_leaf_110_core_clock immu_0.page_table\[12\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3633_ _0812_ net258 _1320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4517__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5714__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4073__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3564_ _1218_ _1281_ _1282_ net533 net542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6352_ _0734_ clknet_leaf_71_core_clock immu_1.page_table\[13\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5303_ _1977_ _2189_ _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_80_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6283_ _0665_ clknet_leaf_34_core_clock dmmu0.page_table\[0\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3495_ net51 dmmu0.long_off_reg\[6\] _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6100__I _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5234_ _2455_ _2470_ _2472_ net1021 _2476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5165_ _2431_ _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4116_ _1770_ _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5096_ _2390_ _0115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6905__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4047_ _1306_ _1696_ _1706_ _1707_ net673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4453__A1 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input211_I core_reset vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input309_I ic0_wb_adr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4205__A1 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5998_ _2917_ _0490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5953__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _2305_ _0053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_1811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6619_ _0192_ clknet_leaf_17_core_clock immu_0.page_table\[0\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6435__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7106__I net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6010__I _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6130__A1 net559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output430_I net430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output528_I net528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4692__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6585__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3878__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4747__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3558__I0 net160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3802__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6121__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3280_ _0948_ _1022_ _1025_ _0875_ _1026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__6928__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4683__A1 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5880__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6970_ _0543_ clknet_leaf_58_core_clock dmmu1.page_table\[0\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4435__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5921_ _1770_ _2872_ _2874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_76_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4986__A2 _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5852_ net94 _2818_ _2820_ dmmu0.page_table\[1\]\[11\] _2833_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6308__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4803_ _2212_ _0000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5935__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5783_ _1863_ _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_72_910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4734_ _1819_ _2157_ _2159_ immu_0.page_table\[15\]\[9\] _2169_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4665_ _2128_ _0755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6458__CLK clknet_leaf_23_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6404_ _0786_ clknet_leaf_106_core_clock immu_0.page_table\[14\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3616_ _1311_ net693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4596_ _2086_ _0728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4371__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6335_ _0717_ clknet_leaf_75_core_clock immu_1.page_table\[15\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3547_ _1273_ net544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input161_I c1_o_mem_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input259_I dcache_wb_o_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6266_ _0648_ clknet_leaf_83_core_clock immu_1.page_table\[4\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3478_ net156 dmmu1.long_off_reg\[6\] _1216_ _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_50_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5217_ _2328_ _2447_ _2449_ net954 _2465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6197_ _0579_ clknet_leaf_1_core_clock immu_0.page_table\[11\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4674__A1 _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5148_ _2421_ _0136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input22_I c0_o_mem_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5079_ _2332_ _2366_ _2368_ net1014 _2380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output478_I net478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_1772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6103__A1 _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_2072 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1934 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5862__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3313__B _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4968__A2 _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1055 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5917__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3539__I _1269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6600__CLK clknet_leaf_17_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4028__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4450_ net95 _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__5145__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold207 dmmu1.page_table\[5\]\[8\] net941 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold218 dmmu0.page_table\[14\]\[2\] net952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6750__CLK clknet_leaf_28_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold229 dmmu0.page_table\[1\]\[2\] net963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4353__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3401_ _1140_ _1122_ _1141_ _1142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_65_1872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4381_ _1866_ _1942_ _1944_ net964 _1953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_1260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3332_ _1072_ _1073_ _1074_ _1075_ _0877_ _0878_ _1076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_6120_ _2986_ _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6051_ _2788_ _2941_ _2943_ dmmu1.page_table\[2\]\[4\] _2948_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3263_ _0899_ dmmu1.page_table\[12\]\[4\] _1009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4656__A1 _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5002_ _2335_ _0076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3194_ _0940_ _0942_ _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4120__A3 _0815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_42_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6953_ _0526_ clknet_leaf_57_core_clock dmmu1.page_table\[1\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5904_ _2864_ _0449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6884_ _0457_ clknet_leaf_48_core_clock dmmu1.page_table\[6\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3631__A2 net257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5835_ _2824_ _0420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6280__CLK clknet_leaf_37_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5766_ _2782_ _2778_ _2780_ dmmu1.page_table\[10\]\[1\] _2783_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5384__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3395__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4717_ _2160_ _0775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5697_ _2741_ _0365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input376_I ic1_wb_adr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4648_ _2069_ _2108_ _2110_ net877 _2118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_2061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_884 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4579_ _2051_ _2075_ _2077_ immu_1.page_table\[14\]\[0\] _2078_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6318_ _0700_ clknet_leaf_70_core_clock dmmu1.page_table\[14\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_1967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_1208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6249_ _0631_ clknet_leaf_88_core_clock immu_1.page_table\[5\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5844__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3870__A2 net238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output595_I net595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6773__CLK clknet_leaf_103_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3386__A1 net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3481__S1 _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6175__I1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3094__I _0849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3233__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3689__A2 net310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_73_2390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4638__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput350 ic1_mem_data[27] net350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput361 ic1_mem_data[8] net361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput372 ic1_wb_adr[3] net372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput383 ic1_wb_we net383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_26_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput394 inner_wb_i_dat[14] net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold90 dmmu0.page_table\[2\]\[3\] net824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3861__A2 _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5063__A1 _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3950_ net112 immu_1.high_addr_off\[2\] _1613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4810__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3613__A2 net263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ _1502_ _1539_ _1545_ _1408_ _1546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_6_1382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5620_ _1976_ _2412_ _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_6_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3377__A1 net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5551_ _2529_ _2647_ _2649_ net998 _2659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4502_ _2026_ _0694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5118__A2 _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5482_ _2620_ _0271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3218__B _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4433_ _1806_ _1979_ _1982_ dmmu0.page_table\[0\]\[4\] _1987_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_6_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3224__S1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7152_ net392 net607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4364_ _1943_ _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6079__B1 _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6103_ _1823_ _2975_ _2977_ dmmu1.page_table\[0\]\[0\] _2978_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3315_ _0938_ _1059_ _1060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_6_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4295_ _1857_ _1894_ _1897_ immu_1.page_table\[0\]\[5\] _1903_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7083_ net336 net489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6034_ _2937_ _0506_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_52_1762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3246_ _0908_ dmmu1.page_table\[4\]\[4\] _0992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_52_1773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3301__A1 _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_2027 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3177_ _0897_ _0925_ _0926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_2038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input124_I c1_o_mem_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Left_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_1_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4563__I _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6936_ _0509_ clknet_leaf_51_core_clock dmmu1.page_table\[2\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6796__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6867_ _0440_ clknet_leaf_65_core_clock dmmu1.page_table\[8\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5818_ _2103_ _2802_ _2804_ net789 _2814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6798_ _0371_ clknet_leaf_49_core_clock dmmu1.page_table\[12\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5749_ _2771_ _0387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4317__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3215__S1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4868__A1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4738__I net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7114__I net390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5293__A1 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output510_I net510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5045__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5596__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5348__A2 _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3359__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3454__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6519__CLK clknet_leaf_109_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_2327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_71_2338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6669__CLK clknet_leaf_104_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5808__B1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3100_ net132 net27 _0850_ _0853_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4080_ _1502_ _1737_ _1739_ _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_78_1348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3031_ _0811_ net559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_69_2267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput180 c1_o_req_ppl_submit net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_1613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput191 c1_sr_bus_addr[4] net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_1624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_2278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3390__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_2044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4982_ _2271_ _2317_ _2319_ dmmu0.page_table\[14\]\[4\] _2324_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5587__A2 _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6721_ _0294_ clknet_leaf_37_core_clock dmmu0.page_table\[3\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3933_ immu_1.page_table\[12\]\[6\] immu_1.page_table\[13\]\[6\] immu_1.page_table\[14\]\[6\]
+ immu_1.page_table\[15\]\[6\] _1474_ _1433_ _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_59_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinterconnect_inner_708 c0_i_core_int_sreg[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_74_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_inner_719 c0_i_core_int_sreg[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_6652_ _0225_ clknet_leaf_24_core_clock dmmu0.page_table\[11\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3864_ immu_0.page_table\[12\]\[4\] immu_0.page_table\[13\]\[4\] immu_0.page_table\[14\]\[4\]
+ immu_0.page_table\[15\]\[4\] _1463_ _1371_ _1530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_73_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5603_ _2689_ _0323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_41_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6583_ _0156_ clknet_leaf_21_core_clock immu_0.page_table\[3\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3795_ _1369_ _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6199__CLK clknet_leaf_2_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5534_ _2650_ _0293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_1775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5465_ immu_1.high_addr_off\[6\] _1861_ _2603_ _2610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput610 net610 ic0_wb_i_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput621 net621 ic1_mem_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput632 net632 ic1_mem_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_41_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4416_ net90 _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
Xoutput643 net643 ic1_wb_i_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5511__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput654 net654 ic1_wb_i_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5396_ net86 _1787_ _1971_ _1972_ _2569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
Xoutput665 net665 inner_wb_adr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_2086 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput676 net676 inner_wb_adr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3522__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7135_ net65 net588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput687 net687 inner_wb_o_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1948 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4347_ _1855_ _1927_ _1929_ immu_1.page_table\[5\]\[4\] _1934_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput698 net698 inner_wb_o_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_35_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input241_I dcache_wb_adr[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input339_I ic1_mem_data[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7066_ net406 net463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4278_ _1872_ _1825_ _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__5275__A1 net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6017_ _2784_ _2924_ _2926_ dmmu1.page_table\[3\]\[2\] _2929_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3229_ dmmu0.page_table\[0\]\[3\] dmmu0.page_table\[1\]\[3\] dmmu0.page_table\[2\]\[3\]
+ dmmu0.page_table\[3\]\[3\] _0950_ _0952_ _0976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_39_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5027__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3411__B _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_26_core_clock clknet_3_2_0_core_clock clknet_leaf_26_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_48_1639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3589__A1 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4786__B1 _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6919_ _0492_ clknet_leaf_59_core_clock dmmu1.page_table\[4\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_1454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4002__A2 _1663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7109__I net400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3436__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5750__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3761__A1 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6811__CLK clknet_leaf_49_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_65_core_clock clknet_3_6_0_core_clock clknet_leaf_65_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6961__CLK clknet_leaf_62_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3816__A2 _1459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1933 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_1370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__A2 _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_2020 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3124__S0 _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_2006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6341__CLK clknet_leaf_71_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4529__B1 _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3547__I _1273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_2514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3201__B1 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3580_ _1290_ net423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3991__B net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3752__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6491__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5250_ _1971_ _2205_ _2484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_27_1770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ net194 net193 net192 _1836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_43_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5181_ _2440_ _0150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4132_ net85 _1778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_21_2081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5257__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4063_ _1378_ _1720_ _1722_ _1723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_30_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__A1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4965_ _2313_ _0061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_43_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6704_ _0277_ clknet_leaf_39_core_clock dmmu0.page_table\[4\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3916_ net6 immu_0.high_addr_off\[1\] _1580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_30_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4896_ _2267_ _2261_ _2263_ net835 _2268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6635_ _0208_ clknet_leaf_12_core_clock dmmu0.page_table\[12\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3847_ net237 _1513_ _1360_ _1514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6834__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input191_I c1_sr_bus_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input289_I ic0_mem_data[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6566_ _0139_ clknet_leaf_18_core_clock immu_0.page_table\[5\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5732__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3778_ _1440_ _1443_ _1444_ _1445_ _1446_ _1447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_28_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5517_ _2463_ _2630_ _2632_ net932 _2640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6497_ _0070_ clknet_leaf_14_core_clock dmmu0.page_table\[14\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5448_ _1895_ net210 _2599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput440 net440 c0_i_req_data[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input52_I c0_o_mem_high_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput451 net451 c0_i_req_data[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput462 net462 c1_disable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6984__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput473 net473 c1_i_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput484 net484 c1_i_req_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3192__I _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5379_ _2560_ _0228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput495 net495 c1_i_req_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7118_ net394 net571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5248__A1 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6214__CLK clknet_leaf_84_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7049_ net285 net436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_29_Right_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_1229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3354__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_2108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6364__CLK clknet_leaf_77_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4759__B1 _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A1 _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5971__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_2037 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3982__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Right_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3409__S1 _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5184__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4931__B1 _2291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5487__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_Right_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6707__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_47_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_2047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6857__CLK clknet_leaf_98_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4750_ _2180_ _0788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_56_Right_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3701_ net313 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_55_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4681_ _2136_ _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6420_ _0802_ clknet_leaf_108_core_clock immu_0.page_table\[12\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3632_ _1319_ net686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5714__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4073__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3725__A1 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _0733_ clknet_leaf_75_core_clock immu_1.page_table\[13\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3563_ _1154_ _1186_ _1231_ _1282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_64_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5302_ _2514_ _0197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6282_ _0664_ clknet_leaf_33_core_clock dmmu0.page_table\[0\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3494_ _1204_ _1218_ _1232_ net532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__6237__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5233_ _2475_ _0167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_65_Right_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5164_ _1980_ _2429_ _2431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4115_ _1769_ _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5095_ _2273_ _2382_ _2384_ net1073 _2390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6387__CLK clknet_leaf_74_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4046_ _1535_ net244 _1707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__A2 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input204_I c1_sr_bus_data_o[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_74_Right_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4205__A2 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5997_ _2794_ _2907_ _2909_ net1058 _2917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4948_ _2267_ _2299_ _2302_ dmmu0.page_table\[7\]\[2\] _2305_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_1413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5953__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3964__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4879_ _2255_ _0033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6618_ _0191_ clknet_leaf_5_core_clock immu_0.page_table\[0\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5166__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6549_ _0122_ clknet_leaf_7_core_clock immu_0.page_table\[6\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4913__B1 _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3915__I net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5469__A1 _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3851__S _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4692__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7122__I net67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3878__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_1701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_4_Left_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_2056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3097__I _0851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5157__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3558__I1 net55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3802__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4683__A2 _2137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5880__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7032__I net277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4435__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A1 _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5920_ _2872_ _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_18_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_3_0_core_clock clknet_0_core_clock clknet_3_3_0_core_clock vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_17_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ _2832_ _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4802_ _1797_ _2208_ _2210_ immu_0.page_table\[13\]\[1\] _2212_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5782_ _2793_ _0398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5935__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3946__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4733_ _2168_ _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4664_ _2059_ _2123_ _2125_ immu_1.page_table\[11\]\[2\] _2128_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6403_ _0785_ clknet_leaf_105_core_clock immu_0.page_table\[15\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3615_ _1308_ net264 _1311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3735__I _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4595_ _1866_ _2075_ _2077_ net752 _2086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_1662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4371__A1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6334_ _0716_ clknet_leaf_61_core_clock immu_1.page_table\[15\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3546_ net135 net30 _1267_ _1273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ _0647_ clknet_leaf_84_core_clock immu_1.page_table\[4\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3477_ _1187_ _1190_ _1215_ _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5950__I _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input154_I c1_o_mem_high_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5216_ _2464_ _0161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6196_ _0578_ clknet_leaf_108_core_clock immu_0.page_table\[11\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4674__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4566__I _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5147_ _2271_ _2414_ _2416_ net1069 _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_2047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input321_I ic0_wb_adr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5078_ _2379_ _0108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input15_I c0_o_mem_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4029_ _1439_ _1689_ _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3937__A1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6402__CLK clknet_leaf_107_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5139__B1 _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7117__I net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6552__CLK clknet_leaf_4_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6103__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_2084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5311__B1 _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5614__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5465__I1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__B1 _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3928__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4028__S1 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3555__I _1277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold208 dmmu1.page_table\[2\]\[1\] net942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold219 immu_0.page_table\[3\]\[7\] net953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4353__A1 _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3400_ net48 dmmu0.long_off_reg\[3\] _1141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_22_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4380_ _1952_ _0646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_885 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3331_ dmmu0.page_table\[8\]\[6\] dmmu0.page_table\[9\]\[6\] dmmu0.page_table\[10\]\[6\]
+ dmmu0.page_table\[11\]\[6\] _0864_ _0941_ _1075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_61_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4105__A1 _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6050_ _2947_ _0512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3262_ dmmu1.page_table\[13\]\[4\] _1008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_1412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I c0_o_instr_long_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4656__A2 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ _1996_ _2316_ _2318_ net995 _2335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3193_ dmmu0.page_table\[4\]\[1\] dmmu0.page_table\[5\]\[1\] dmmu0.page_table\[6\]\[1\]
+ dmmu0.page_table\[7\]\[1\] _0864_ _0941_ _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_79_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ _0525_ clknet_leaf_52_core_clock dmmu1.page_table\[1\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_2086 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5903_ _2790_ _2856_ _2858_ dmmu1.page_table\[7\]\[5\] _2864_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6883_ _0456_ clknet_leaf_66_core_clock dmmu1.page_table\[7\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6425__CLK clknet_leaf_105_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5834_ _1799_ _2819_ _2821_ net963 _2824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5765_ _1845_ _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_8_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4716_ _1777_ _2157_ _2159_ immu_0.page_table\[15\]\[0\] _2160_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3395__A2 _1131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5696_ _2049_ _2725_ _2727_ net1043 _2741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6575__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4647_ _2117_ _0748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_2002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3465__I _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input271_I dcache_wb_o_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5541__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input369_I ic1_wb_adr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4578_ _2076_ _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_40_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_2079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6317_ _0699_ clknet_leaf_96_core_clock dmmu1.page_table\[14\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3529_ net142 net37 _0850_ _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6097__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6248_ _0630_ clknet_leaf_88_core_clock immu_1.page_table\[5\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5844__A1 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6179_ dmmu1.long_off_reg\[4\] _1855_ _3016_ _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_2006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6021__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output490_I net490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6918__CLK clknet_leaf_59_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output588_I net588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4583__A1 _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4335__A1 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5590__I _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_1456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4638__A2 _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput340 ic1_mem_data[18] net340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3846__B1 _1503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput351 ic1_mem_data[28] net351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput362 ic1_mem_data[9] net362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput373 ic1_wb_adr[4] net373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xhold80 dmmu0.page_table\[2\]\[7\] net814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput384 inner_disable net384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput395 inner_wb_i_dat[15] net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold91 immu_1.page_table\[10\]\[2\] net825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6448__CLK clknet_leaf_10_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5063__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3074__A1 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4271__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4810__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3880_ _1502_ _1542_ _1544_ _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_39_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6598__CLK clknet_leaf_16_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5765__I _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5550_ _2658_ _0301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4501_ _1868_ _2014_ _2016_ net845 _2026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5481_ _2457_ _2613_ _2615_ dmmu0.page_table\[4\]\[4\] _2620_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4432_ _1986_ _0664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5523__B1 _2631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7151_ net391 net606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4363_ _1912_ _1941_ _1943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6079__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6102_ _2976_ _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3314_ dmmu0.page_table\[4\]\[5\] dmmu0.page_table\[5\]\[5\] dmmu0.page_table\[6\]\[5\]
+ dmmu0.page_table\[7\]\[5\] _0872_ _0941_ _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_10_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7082_ net335 net488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4294_ _1902_ _0610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5826__A1 _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6033_ _2851_ _2923_ _2925_ net858 _2937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3245_ dmmu1.page_table\[5\]\[4\] _0991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_52_1763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3176_ dmmu1.page_table\[4\]\[1\] dmmu1.page_table\[5\]\[1\] dmmu1.page_table\[6\]\[1\]
+ dmmu1.page_table\[7\]\[1\] _0908_ _0910_ _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_33_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_16_core_clock clknet_3_0_0_core_clock clknet_leaf_16_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_1_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input117_I c1_o_instr_long_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6935_ _0508_ clknet_leaf_63_core_clock dmmu1.page_table\[3\]\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6866_ _0439_ clknet_leaf_65_core_clock dmmu1.page_table\[8\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6003__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5817_ _2813_ _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_1079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6797_ _0370_ clknet_leaf_44_core_clock dmmu1.page_table\[12\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_903 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5748_ _2101_ _2760_ _2762_ dmmu1.page_table\[11\]\[8\] _2771_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input82_I c0_sr_bus_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5679_ _2732_ _0356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_66_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_969 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4317__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4868__A2 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_55_core_clock clknet_3_7_0_core_clock clknet_leaf_55_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_77_1530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5293__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output503_I net503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3798__C _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7130__I net60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5045__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3359__A2 _1101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__CLK clknet_leaf_54_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_94_core_clock clknet_3_4_0_core_clock clknet_leaf_94_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_1665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4308__A1 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5505__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_2453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_2464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5808__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6270__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3030_ _0809_ _0810_ mem_dcache_arb.transfer_active _0811_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput170 c1_o_req_addr[15] net170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput181 c1_sr_bus_addr[0] net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_69_2268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput192 c1_sr_bus_addr[5] net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7040__I net307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3390__S1 _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_104_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3047__A1 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4981_ _2323_ _0067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3932_ _1440_ _1595_ _1596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6720_ _0293_ clknet_leaf_34_core_clock dmmu0.page_table\[3\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_1967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6651_ _0224_ clknet_leaf_27_core_clock dmmu0.page_table\[11\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinterconnect_inner_709 c0_i_core_int_sreg[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_3863_ _1368_ _1528_ _1529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5602_ _2457_ _2681_ _2684_ dmmu0.page_table\[6\]\[4\] _2689_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_1691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6582_ _0155_ clknet_leaf_5_core_clock immu_0.page_table\[3\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_41_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5744__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3794_ _1385_ immu_0.page_table\[14\]\[2\] _1462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5533_ _2444_ _2647_ _2649_ net842 _2650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5464_ _2609_ _0264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput600 net600 ic0_mem_req vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_44_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput611 net611 ic0_wb_i_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput622 net622 ic1_mem_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_58_1950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4415_ _1971_ _1972_ _1973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xoutput633 net633 ic1_mem_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_54_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5395_ _2568_ _0236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput644 net644 ic1_wb_i_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_54_1814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6613__CLK clknet_leaf_9_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput655 net655 ic1_wb_i_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput666 net666 inner_wb_adr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7134_ net64 net587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput677 net677 inner_wb_adr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1987 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4346_ _1933_ _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput688 net688 inner_wb_o_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput699 net699 inner_wb_o_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7065_ net211 net461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4277_ _1823_ _1890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input234_I dcache_wb_adr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6016_ _2928_ _0497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3228_ dmmu0.page_table\[4\]\[3\] dmmu0.page_table\[5\]\[3\] dmmu0.page_table\[6\]\[3\]
+ dmmu0.page_table\[7\]\[3\] _0950_ _0952_ _0975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_20_1061 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6763__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4483__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3159_ _0900_ _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_68_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input401_I inner_wb_i_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3038__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4786__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3589__A2 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6918_ _0491_ clknet_leaf_59_core_clock dmmu1.page_table\[4\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5983__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6849_ _0422_ clknet_leaf_34_core_clock dmmu0.page_table\[1\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwire705 _1407_ net705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_52_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3854__S _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3761__A2 _1429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output453_I net453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6293__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7125__I net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4710__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3816__A3 _1468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_2121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_2132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3124__S1 _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_2018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4529__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_2504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3201__B2 _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6636__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6151__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4200_ net191 _1835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_1624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5180_ _2277_ _2430_ _2432_ net852 _2440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6786__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_79_Left_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4131_ _1776_ _1777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_21_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5257__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4062_ _1366_ _1721_ _1722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_1370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4465__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_939 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4217__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5965__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4964_ _1821_ _2298_ _2301_ dmmu0.page_table\[7\]\[10\] _2313_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6703_ _0276_ clknet_leaf_39_core_clock dmmu0.page_table\[4\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3915_ net2 _1579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_19_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4895_ _1799_ _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3440__A1 net50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3846_ _1422_ _1490_ _1498_ _1503_ _1512_ _1513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6634_ _0207_ clknet_leaf_13_core_clock dmmu0.page_table\[12\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_880 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3777_ _1415_ _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_6565_ _0138_ clknet_leaf_20_core_clock immu_0.page_table\[5\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input184_I c1_sr_bus_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5516_ _2639_ _0286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6496_ _0069_ clknet_leaf_24_core_clock dmmu0.page_table\[14\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5447_ net325 _1766_ _2598_ _1771_ _0258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput430 net430 c0_i_req_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_37_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput441 net441 c0_i_req_data[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input351_I ic1_mem_data[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput452 net452 c0_i_req_data[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput463 net463 c1_i_core_int_sreg[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5378_ _2457_ _2553_ _2555_ dmmu0.page_table\[11\]\[4\] _2560_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput474 net474 c1_i_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput485 net485 c1_i_req_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input45_I c0_o_mem_high_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput496 net496 c1_i_req_data[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_6_core_clock clknet_3_0_0_core_clock clknet_leaf_6_core_clock vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7117_ net393 net570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4329_ _1866_ _1911_ _1914_ net1029 _1923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_22_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5248__A2 _2469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7048_ net284 net435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3354__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6509__CLK clknet_leaf_109_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4759__A1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_102_core_clock clknet_3_1_0_core_clock clknet_leaf_102_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5420__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6659__CLK clknet_leaf_23_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5708__B1 _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3982__A2 _1639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5184__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__A1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4931__B2 _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5487__A2 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3498__A1 net52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3670__A1 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_2015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3700_ _1369_ _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_71_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ _2105_ _2122_ _2124_ immu_1.page_table\[11\]\[10\] _2136_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_50_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _0812_ net257 _1319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_1194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6350_ _0732_ clknet_leaf_61_core_clock immu_1.page_table\[13\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3562_ _1169_ _1202_ _1281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5301_ net93 _2501_ _2503_ immu_0.page_table\[0\]\[10\] _2514_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_3_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6281_ _0663_ clknet_leaf_36_core_clock dmmu0.page_table\[0\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3493_ _1219_ _1231_ _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5232_ _2453_ _2470_ _2472_ immu_0.page_table\[2\]\[2\] _2475_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3489__A1 net50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5163_ _2429_ _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4114_ net211 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5094_ _2389_ _0114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4045_ net2 _1700_ _1705_ _1382_ _1422_ _1706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__4453__A3 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3661__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6801__CLK clknet_leaf_42_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5996_ _2916_ _0489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4947_ _2304_ _0052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input399_I inner_wb_i_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3964__A2 _1626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4878_ _1821_ _2241_ _2243_ net745 _2255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5166__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6617_ _0190_ clknet_leaf_15_core_clock immu_0.page_table\[0\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3829_ _1372_ _1492_ _1495_ _1366_ _1496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_43_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4913__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6548_ _0121_ clknet_leaf_3_core_clock immu_0.page_table\[6\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1966 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6115__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6479_ _0052_ clknet_leaf_32_core_clock dmmu0.page_table\[7\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6331__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4429__B1 _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_2031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1016 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_1303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3652__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6481__CLK clknet_leaf_29_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__B1 _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_2092 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5157__A1 _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_1_0_core_clock_I clknet_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4668__B1 _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5880__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6824__CLK clknet_leaf_48_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5093__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3643__A1 _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_909 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5768__I _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5850_ _2531_ _2818_ _2820_ net1034 _2832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4801_ _2211_ _0808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5396__A1 net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6974__CLK clknet_leaf_62_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5781_ _2792_ _2778_ _2780_ net763 _2793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4732_ _1817_ _2157_ _2159_ net919 _2168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3946__A2 _1605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4663_ _2127_ _0754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6204__CLK clknet_leaf_93_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6402_ _0784_ clknet_leaf_107_core_clock immu_0.page_table\[15\]\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3614_ _1310_ net692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_883 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4594_ _2085_ _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3237__B _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3545_ _1272_ net558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4371__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6333_ _0715_ clknet_leaf_71_core_clock immu_1.page_table\[15\]\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6264_ _0646_ clknet_leaf_84_core_clock immu_1.page_table\[4\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3476_ net155 dmmu1.long_off_reg\[5\] _1215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6354__CLK clknet_leaf_75_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5215_ _2463_ _2447_ _2449_ net953 _2464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6195_ _0577_ clknet_leaf_109_core_clock immu_0.page_table\[11\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input147_I c1_o_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5146_ _2420_ _0135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3882__A1 net110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5077_ _2330_ _2367_ _2369_ net860 _2379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input314_I ic0_wb_adr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4028_ immu_1.page_table\[8\]\[9\] immu_1.page_table\[9\]\[9\] immu_1.page_table\[10\]\[9\]
+ immu_1.page_table\[11\]\[9\] _1409_ _1410_ _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_75_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1000 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4831__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ _1873_ _1892_ _2030_ _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_48_986 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5139__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_2019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_894 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_2090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output533_I net533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5311__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7133__I net63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6847__CLK clknet_leaf_36_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5075__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5614__A2 _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3625__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6997__CLK clknet_leaf_95_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3102__S _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5378__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_109_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6227__CLK clknet_leaf_87_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_975 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4050__A1 net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6377__CLK clknet_leaf_73_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold209 immu_1.page_table\[15\]\[4\] net943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_65_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4353__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3330_ dmmu0.page_table\[12\]\[6\] dmmu0.page_table\[13\]\[6\] dmmu0.page_table\[14\]\[6\]
+ dmmu0.page_table\[15\]\[6\] _0864_ _0941_ _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_1_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4105__A2 net381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3261_ _0889_ _1005_ _1006_ _1007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7043__I net279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_59_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5000_ _2334_ _0075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4656__A3 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3192_ _0867_ _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_79_1060 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6951_ _0524_ clknet_leaf_51_core_clock dmmu1.page_table\[1\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5902_ _2863_ _0448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6882_ _0455_ clknet_leaf_65_core_clock dmmu1.page_table\[7\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5833_ _2823_ _0419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_1075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5764_ _2781_ _0392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_956 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4715_ _2158_ _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5695_ _2740_ _0364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4646_ _2067_ _2108_ _2110_ net929 _2117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5541__A1 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4577_ _1912_ _2074_ _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_1340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input264_I dcache_wb_o_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6316_ _0698_ clknet_leaf_69_core_clock dmmu1.page_table\[14\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3528_ _1263_ net550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_45_core_clock clknet_3_6_0_core_clock clknet_leaf_45_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6097__A2 _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6247_ _0629_ clknet_leaf_84_core_clock immu_1.page_table\[5\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3459_ _0906_ _1198_ _1199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_1070 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5844__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6178_ _3020_ _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_24_Left_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5129_ _2409_ _0129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5402__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_2001 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4804__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_2089 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A1 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_61_core_clock_I clknet_3_7_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6021__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4032__A1 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3466__S0 _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_33_Left_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4583__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7128__I net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_84_core_clock clknet_3_5_0_core_clock clknet_leaf_84_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4335__A2 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_73_2392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4099__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_42_Left_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput330 ic1_mem_ack net330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3846__A1 _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput341 ic1_mem_data[19] net341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput352 ic1_mem_data[29] net352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_1777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput363 ic1_wb_adr[0] net363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput374 ic1_wb_adr[5] net374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_1807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput385 inner_embed_mode net385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xhold70 dmmu1.page_table\[2\]\[12\] net804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold81 immu_0.page_table\[14\]\[10\] net815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput396 inner_wb_i_dat[1] net396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold92 immu_1.page_table\[15\]\[5\] net826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_37_1206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4271__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3074__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Left_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7038__I net305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4500_ _2025_ _0693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5480_ _2619_ _0270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3209__S0 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_1 net383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4431_ _1803_ _1979_ _1982_ dmmu0.page_table\[0\]\[3\] _1986_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5523__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4362_ _1941_ _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_26_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7150_ net390 net605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6079__A2 _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6101_ _1770_ _2974_ _2976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_60_Left_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3313_ _0940_ _1057_ _0958_ _1058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7081_ net334 net487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4293_ _1854_ _1894_ _1897_ immu_1.page_table\[0\]\[4\] _1902_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_24_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5287__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6032_ _2936_ _0505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3244_ dmmu1.page_table\[6\]\[4\] dmmu1.page_table\[7\]\[4\] _0908_ _0990_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_52_1764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3175_ _0922_ _0923_ _0907_ _0924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_2018 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5039__B1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_2029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6934_ _0507_ clknet_leaf_57_core_clock dmmu1.page_table\[3\]\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4065__C _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6542__CLK clknet_leaf_19_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6865_ _0438_ clknet_leaf_42_core_clock dmmu1.page_table\[8\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6003__A2 _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5816_ _2101_ _2802_ _2804_ dmmu1.page_table\[9\]\[8\] _2813_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4014__A1 _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6796_ _0369_ clknet_leaf_45_core_clock dmmu1.page_table\[12\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5747_ _2770_ _0386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input381_I ic1_wb_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6692__CLK clknet_leaf_91_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5678_ _2061_ _2726_ _2728_ dmmu1.page_table\[13\]\[3\] _2732_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input75_I c0_o_req_ppl_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4317__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ _2106_ _0741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_66_1479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1029 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3828__A1 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1936 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4253__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4005__A1 net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6190__C _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_2590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5505__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4308__A2 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_2454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1953 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6415__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__B1 _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5808__A2 _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput160 c1_o_mem_sel[0] net160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3295__A2 _1040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput171 c1_o_req_addr[1] net171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput182 c1_sr_bus_addr[10] net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_1615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_2269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput193 c1_sr_bus_addr[6] net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6565__CLK clknet_leaf_20_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_2024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _2269_ _2317_ _2319_ net926 _2323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3047__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3931_ immu_1.page_table\[8\]\[6\] immu_1.page_table\[9\]\[6\] immu_1.page_table\[10\]\[6\]
+ immu_1.page_table\[11\]\[6\] _1474_ _1433_ _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_74_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6650_ _0223_ clknet_leaf_10_core_clock dmmu0.page_table\[15\]\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3862_ immu_0.page_table\[8\]\[4\] immu_0.page_table\[9\]\[4\] immu_0.page_table\[10\]\[4\]
+ immu_0.page_table\[11\]\[4\] _1463_ _1391_ _1528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_58_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5601_ _2688_ _0322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5744__A1 _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ _0154_ clknet_leaf_4_core_clock immu_0.page_table\[3\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_41_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3793_ immu_0.page_table\[12\]\[2\] immu_0.page_table\[13\]\[2\] _1396_ _1461_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5532_ _2648_ _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_14_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3850__S0 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5463_ immu_1.high_addr_off\[5\] _1858_ _2603_ _2609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput601 net601 ic0_rst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_58_1940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput612 net612 ic0_wb_i_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_48_1198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4414_ net83 net76 _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_26_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput623 net623 ic1_mem_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput634 net634 ic1_mem_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5394_ _1996_ _2552_ _2554_ dmmu0.page_table\[11\]\[12\] _2568_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput645 net645 ic1_wb_i_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_22_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_1906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput656 net656 ic1_wb_i_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_54_1815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7133_ net63 net586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput667 net667 inner_wb_adr[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4180__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4345_ _1852_ _1927_ _1929_ net1085 _1933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput678 net678 inner_wb_adr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput689 net689 inner_wb_o_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_35_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4276_ _1889_ _0605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7064_ net276 net460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_35_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6908__CLK clknet_leaf_64_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _2782_ _2924_ _2926_ dmmu1.page_table\[3\]\[1\] _2928_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3227_ _0883_ _0973_ _0879_ _0974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4855__I _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4483__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5680__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input227_I dcache_mem_o_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3158_ _0898_ _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3038__A2 _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3089_ net127 net22 _0842_ _0847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5432__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6917_ _0490_ clknet_leaf_55_core_clock dmmu1.page_table\[4\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5983__A1 _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4786__A2 _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6848_ _0421_ clknet_leaf_45_core_clock dmmu0.page_table\[1\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1899 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6779_ _0352_ clknet_leaf_99_core_clock dmmu0.long_off_reg\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_21_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_2106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output446_I net446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4710__A2 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6588__CLK clknet_leaf_14_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7141__I net396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_2122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3029__A2 net159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_2008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4529__A2 _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5726__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_2505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_2527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3832__S0 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6151__A1 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3780__S _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4130_ net92 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_20_995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_2083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4061_ immu_0.page_table\[12\]\[10\] immu_0.page_table\[13\]\[10\] immu_0.page_table\[14\]\[10\]
+ immu_0.page_table\[15\]\[10\] _1487_ _1390_ _1721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_30_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7051__I net287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4465__A1 _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1994 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4217__A1 _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5965__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4963_ _2312_ _0060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6702_ _0275_ clknet_leaf_45_core_clock dmmu0.page_table\[4\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_1129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3914_ net659 _1577_ _1578_ net668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_28_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4894_ _2266_ _0037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_15_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6633_ _0206_ clknet_leaf_23_core_clock dmmu0.page_table\[12\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3845_ _0813_ _1511_ _1512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4076__S0 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6564_ _0137_ clknet_leaf_20_core_clock immu_0.page_table\[5\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3776_ immu_1.page_table\[2\]\[1\] immu_1.page_table\[3\]\[1\] _1435_ _1445_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5515_ _2461_ _2630_ _2632_ net1087 _2639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_873 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6495_ _0068_ clknet_leaf_29_core_clock dmmu0.page_table\[14\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input177_I c1_o_req_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5446_ _1422_ net379 _2598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput420 net420 c0_i_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_37_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput431 net431 c0_i_req_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput442 net442 c0_i_req_data[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6730__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput453 net453 c0_i_req_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4153__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput464 net464 c1_i_core_int_sreg[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput475 net475 c1_i_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_1102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5377_ _2559_ _0227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input344_I ic1_mem_data[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput486 net486 c1_i_req_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7116_ net392 net569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput497 net497 c1_i_req_data[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4328_ _1922_ _0624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input38_I c0_o_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ net283 net434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4259_ _1849_ _1876_ _1878_ net983 _1881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_57_1209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5410__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_2090 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4759__A2 _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1952 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_2039 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5708__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6260__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5184__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output563_I net563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4931__A2 _2290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1024 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6040__I _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6133__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3670__A2 net321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1006 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5947__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1954 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6603__CLK clknet_leaf_5_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3630_ _1318_ net700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3186__A1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6753__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3561_ _1280_ net561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7046__I net282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ _2513_ _0196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1015 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1878 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3507__C _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3492_ _0883_ _1223_ _1227_ _1230_ _1119_ _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_6280_ _0662_ clknet_leaf_37_core_clock dmmu0.page_table\[0\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_1168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5231_ _2474_ _0166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4686__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5162_ _1789_ _2428_ _2429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4113_ net659 _1767_ _1768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5093_ _2271_ _2382_ _2384_ immu_0.page_table\[7\]\[4\] _2389_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4044_ _1701_ _1702_ _1703_ _1704_ _1367_ _1383_ _1705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_79_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3110__A1 net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3661__A2 net373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5995_ _2792_ _2907_ _2909_ net977 _2916_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6283__CLK clknet_leaf_34_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4946_ _2265_ _2299_ _2302_ dmmu0.page_table\[7\]\[1\] _2304_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3413__A2 _1153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_66_core_clock_I clknet_3_6_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4877_ _2254_ _0032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_1836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input294_I ic0_mem_data[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6616_ _0189_ clknet_leaf_15_core_clock immu_0.page_table\[0\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3828_ _1391_ _1493_ _1494_ _1495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5166__A2 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3177__A1 _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6547_ _0120_ clknet_leaf_8_core_clock immu_0.page_table\[7\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3759_ immu_0.page_table\[6\]\[1\] immu_0.page_table\[7\]\[1\] immu_0.page_table\[14\]\[1\]
+ immu_0.page_table\[15\]\[1\] _1370_ _1377_ _1428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__4913__A2 _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6115__A1 _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6478_ _0051_ clknet_leaf_27_core_clock dmmu0.page_table\[7\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5429_ _2589_ _0249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_7_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5874__B1 _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4429__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5626__B1 _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6626__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3652__A2 net371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A1 _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6051__B1 _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_932 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4601__A1 _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output680_I net680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6776__CLK clknet_leaf_100_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_998 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5157__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4365__B1 _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_929 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3327__C _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4668__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3340__A1 net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5093__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3643__A2 net363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _1777_ _2208_ _2210_ net1016 _2211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5780_ _1860_ _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_8_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_965 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4731_ _2167_ _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4662_ _2057_ _2123_ _2125_ immu_1.page_table\[11\]\[1\] _2127_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6401_ _0783_ clknet_leaf_107_core_clock immu_0.page_table\[15\]\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3613_ _1308_ net263 _1310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _2069_ _2075_ _2077_ net1007 _2085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_1511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6332_ _0714_ clknet_leaf_75_core_clock immu_1.page_table\[15\]\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3544_ net149 net44 _1267_ _1272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_35_core_clock clknet_3_3_0_core_clock clknet_leaf_35_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6263_ _0645_ clknet_leaf_86_core_clock immu_1.page_table\[4\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3475_ _1211_ _1213_ _0895_ _1214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_0_951 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5214_ _1814_ _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6194_ _0576_ clknet_leaf_8_core_clock immu_0.page_table\[11\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5145_ _2269_ _2414_ _2416_ immu_0.page_table\[5\]\[3\] _2420_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6649__CLK clknet_leaf_12_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5608__B1 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5076_ _2378_ _0107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4027_ _1686_ _1687_ _1416_ _1688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4831__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input307_I ic0_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6799__CLK clknet_leaf_50_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5978_ _2905_ _0482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3398__A1 _1118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4595__B1 _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4929_ _1788_ _2240_ _2284_ _2290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_62_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_74_core_clock clknet_3_5_0_core_clock clknet_leaf_74_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5139__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4347__B1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3428__B _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1931 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5311__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1926 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3163__B _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output526_I net526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5075__A1 _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3625__A2 net269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1025 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5378__A2 _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5109__I _2397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1875 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5838__B1 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3260_ _0899_ dmmu1.page_table\[14\]\[4\] _0910_ _1006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3313__A1 _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3191_ _0875_ _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6941__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6950_ _0523_ clknet_leaf_53_core_clock dmmu1.page_table\[1\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5901_ _2788_ _2856_ _2858_ dmmu1.page_table\[7\]\[4\] _2863_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_2077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6881_ _0454_ clknet_leaf_66_core_clock dmmu1.page_table\[7\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6015__B1 _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1988 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5832_ _1796_ _2819_ _2821_ dmmu0.page_table\[1\]\[1\] _2823_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_1398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1043 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5763_ _2776_ _2778_ _2780_ net981 _2781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_1592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4714_ _2140_ _2156_ _2158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5447__C _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5694_ _2047_ _2725_ _2727_ net897 _2740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6321__CLK clknet_leaf_96_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4329__B1 _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4645_ _2116_ _0747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_2026 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4576_ _2074_ _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5541__A2 _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_2048 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_876 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6315_ _0697_ clknet_leaf_70_core_clock dmmu1.page_table\[14\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3527_ net141 net36 _0850_ _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_898 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6471__CLK clknet_leaf_22_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input257_I dcache_wb_o_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6246_ _0628_ clknet_leaf_82_core_clock immu_1.page_table\[5\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3458_ dmmu1.page_table\[8\]\[10\] dmmu1.page_table\[9\]\[10\] dmmu1.page_table\[10\]\[10\]
+ dmmu1.page_table\[11\]\[10\] _0887_ _0900_ _1198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3304__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4501__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6177_ dmmu1.long_off_reg\[3\] _1852_ _3016_ _3020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3389_ _1129_ _1130_ _0896_ _1131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5128_ _2328_ _2398_ _2400_ immu_0.page_table\[6\]\[8\] _2409_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input20_I c0_o_mem_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5057__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5059_ _2258_ _2367_ _2369_ net978 _2370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4804__A1 _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_1432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A2 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1886 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3466__S1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3091__I0 net128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3791__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_916 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6814__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4335__A3 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7144__I net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4099__A2 net275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6964__CLK clknet_leaf_56_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput320 ic0_wb_adr[5] net320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput331 ic1_mem_data[0] net331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3846__A2 _1490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput342 ic1_mem_data[1] net342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput353 ic1_mem_data[2] net353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold60 immu_1.page_table\[2\]\[5\] net794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput364 ic1_wb_adr[10] net364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold71 immu_0.page_table\[12\]\[4\] net805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput375 ic1_wb_adr[6] net375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold82 dmmu0.page_table\[12\]\[2\] net816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput386 inner_ext_irq net386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput397 inner_wb_i_dat[2] net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold93 dmmu0.page_table\[15\]\[10\] net827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_3_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_2042 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4271__A2 _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6344__CLK clknet_leaf_71_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_935 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3782__A1 net705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6494__CLK clknet_leaf_27_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3209__S1 _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4430_ _1985_ _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_2 net383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__A2 _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4361_ _1839_ _1873_ _1892_ _1941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6100_ _2974_ _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3312_ dmmu0.page_table\[0\]\[5\] dmmu0.page_table\[1\]\[5\] dmmu0.page_table\[2\]\[5\]
+ dmmu0.page_table\[3\]\[5\] _0864_ _0941_ _1057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_7080_ net333 net486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4292_ _1901_ _0609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5287__A1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ _2849_ _2924_ _2926_ net780 _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3243_ _0932_ _0892_ _0933_ _0989_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_20_1222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1009 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3174_ dmmu1.page_table\[8\]\[1\] dmmu1.page_table\[9\]\[1\] dmmu1.page_table\[10\]\[1\]
+ dmmu1.page_table\[11\]\[1\] _0908_ _0910_ _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5039__A1 _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6933_ _0506_ clknet_leaf_63_core_clock dmmu1.page_table\[3\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _0437_ clknet_leaf_50_core_clock dmmu1.page_table\[8\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5815_ _2812_ _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6795_ _0368_ clknet_leaf_45_core_clock dmmu1.page_table\[12\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6837__CLK clknet_leaf_48_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1985 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5746_ _2069_ _2760_ _2762_ dmmu1.page_table\[11\]\[7\] _2770_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_1947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4081__C _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1958 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5677_ _2731_ _0355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input374_I ic1_wb_adr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4628_ _2105_ _2089_ _2091_ net1060 _2106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6987__CLK clknet_leaf_79_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input68_I c0_o_req_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4722__B1 _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ _2064_ _0713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5278__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6229_ _0611_ clknet_leaf_86_core_clock immu_1.page_table\[0\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6217__CLK clknet_leaf_83_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_1418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6367__CLK clknet_leaf_61_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1959 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5450__A1 _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_879 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output593_I net593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_2061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7139__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5882__I net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_2591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5505__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4308__A3 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_2444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3335__C _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__A1 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput150 c1_o_mem_high_addr[0] net150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_1575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput161 c1_o_mem_sel[1] net161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput172 c1_o_req_addr[2] net172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3351__B _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput183 c1_sr_bus_addr[11] net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput194 c1_sr_bus_addr[7] net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3930_ _1579_ _1582_ _1593_ _1348_ _1594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3861_ _1375_ _1526_ _1378_ _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7049__I net285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5600_ _2455_ _2681_ _2684_ dmmu0.page_table\[6\]\[3\] _2688_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6580_ _0153_ clknet_leaf_9_core_clock immu_0.page_table\[4\]\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3792_ immu_0.page_table\[4\]\[2\] immu_0.page_table\[5\]\[2\] immu_0.page_table\[6\]\[2\]
+ immu_0.page_table\[7\]\[2\] _1370_ _1372_ _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_41_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5744__A2 _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5531_ _2300_ _2646_ _2648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4952__B1 _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3850__S1 _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5462_ _2608_ _0263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_1729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_2023 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput602 net602 ic0_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3507__A1 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1019 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4413_ net85 net84 _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xoutput613 net613 ic0_wb_i_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4704__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput624 net624 ic1_mem_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5393_ _2567_ _0235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_58_1963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput635 net635 ic1_mem_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput646 net646 ic1_wb_i_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7132_ net62 net585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4180__A1 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput657 net657 ic1_wb_i_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_54_1816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4344_ _1932_ _0630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput668 net668 inner_wb_adr[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput679 net679 inner_wb_adr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7063_ net301 net452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_35_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4275_ _1870_ _1875_ _1877_ immu_1.page_table\[7\]\[10\] _1889_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_35_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6014_ _2927_ _0496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3226_ _0971_ _0972_ _0940_ _0973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4483__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5680__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3157_ _0906_ _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_59_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input122_I c1_o_mem_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3088_ _0846_ net534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3038__A3 _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5432__A1 _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6916_ _0489_ clknet_leaf_54_core_clock dmmu1.page_table\[4\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5983__A2 _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6847_ _0420_ clknet_leaf_36_core_clock dmmu0.page_table\[1\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6778_ _0351_ clknet_leaf_99_core_clock dmmu0.long_off_reg\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_21_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5729_ _2759_ _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_17_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5408__S _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5499__A1 _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_73_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5120__B1 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2003 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_2047 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_2058 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_2123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2012 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_1644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_2009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3985__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3737__A1 net385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_2517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_2528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3832__S1 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6151__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1041 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6532__CLK clknet_leaf_1_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_2062 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_2073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4060_ _1368_ _1719_ _1720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4465__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_908 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4217__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4962_ _1819_ _2299_ _2302_ dmmu0.page_table\[7\]\[9\] _2312_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5965__A2 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6701_ _0274_ clknet_leaf_31_core_clock dmmu0.page_table\[4\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3913_ net659 net239 _1578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_28_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4893_ _2265_ _2261_ _2263_ dmmu0.page_table\[8\]\[1\] _2266_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6632_ _0205_ clknet_leaf_29_core_clock dmmu0.page_table\[12\]\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_15_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5178__B1 _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3844_ _1502_ net705 _1505_ _1510_ _1511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_46_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4076__S1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3728__A1 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_979 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6563_ _0136_ clknet_leaf_18_core_clock immu_0.page_table\[5\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3775_ _1433_ _1439_ _1444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_1531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5514_ _2638_ _0285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6494_ _0067_ clknet_leaf_27_core_clock dmmu0.page_table\[14\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5445_ _2597_ _0257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_1439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput410 net410 c0_i_mem_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_930 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput421 net421 c0_i_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput432 net432 c0_i_req_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput443 net443 c0_i_req_data[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4153__A1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5350__B1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput454 net454 c0_i_req_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5376_ _2455_ _2553_ _2555_ dmmu0.page_table\[11\]\[3\] _2559_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput465 net465 c1_i_mc_core_int vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput476 net476 c1_i_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7115_ net391 net568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput487 net487 c1_i_req_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4327_ _1864_ _1911_ _1914_ net895 _1922_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput498 net498 c1_i_req_data[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3770__I _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input337_I ic1_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7046_ net282 net433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4258_ _1880_ _0596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_1600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3209_ dmmu0.page_table\[0\]\[2\] dmmu0.page_table\[1\]\[2\] dmmu0.page_table\[2\]\[2\]
+ dmmu0.page_table\[3\]\[2\] _0950_ _0952_ _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4189_ _1823_ _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_78_1693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3211__S _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3967__A1 net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5708__A2 _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3719__A1 _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6555__CLK clknet_leaf_18_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_1014 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_896 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_2051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1995 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold190 dmmu1.page_table\[1\]\[11\] net924 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_44_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7152__I net392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5644__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_16_Right_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1034 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_963 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5947__A2 _2872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3502__S0 _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_1977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_905 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3186__A2 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3560_ net161 net56 _0841_ _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_25_Right_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_25_core_clock clknet_3_2_0_core_clock clknet_leaf_25_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_1294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3491_ net51 dmmu0.long_off_reg\[6\] _1229_ _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_51_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5230_ _2451_ _2470_ _2472_ immu_0.page_table\[2\]\[1\] _2474_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5883__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5161_ _1972_ _2296_ _2428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_23_1456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4112_ _1765_ _1766_ _1767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5092_ _2388_ _0113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4043_ immu_0.page_table\[0\]\[9\] immu_0.page_table\[1\]\[9\] immu_0.page_table\[2\]\[9\]
+ immu_0.page_table\[3\]\[9\] _1396_ _1371_ _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_79_1980 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_34_Right_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3741__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6428__CLK clknet_leaf_106_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5994_ _2915_ _0488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_900 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4945_ _2303_ _0051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_23_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4876_ _1819_ _2242_ _2244_ dmmu0.page_table\[9\]\[9\] _2254_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_64_core_clock clknet_3_7_0_core_clock clknet_leaf_64_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_1449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6578__CLK clknet_leaf_18_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3827_ _1463_ immu_0.page_table\[15\]\[3\] _1494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6615_ _0188_ clknet_leaf_6_core_clock immu_0.page_table\[0\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3765__I _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_893 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_Right_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5410__I1 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3177__A2 _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input287_I ic0_mem_data[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6546_ _0119_ clknet_leaf_3_core_clock immu_0.page_table\[7\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3758_ _1382_ _1426_ _1372_ _1427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__5571__B1 _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6477_ _0050_ clknet_leaf_90_core_clock net407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5980__I _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6115__A2 _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3689_ _1350_ net310 _1360_ _1361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_982 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4126__A1 net659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5428_ _2457_ _2582_ _2584_ dmmu0.page_table\[2\]\[4\] _2589_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input50_I c0_o_mem_high_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5874__A1 _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5359_ _2548_ _0220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3206__S _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Right_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5626__A1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4429__A2 _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7029_ net384 net405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_57_1007 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_2099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6051__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4601__A2 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_977 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1073 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_2050 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_61_Right_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_1483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3675__I _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7147__I net402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4365__A1 _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4668__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_70_Right_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_1191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1033 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5093__A2 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6720__CLK clknet_leaf_34_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5396__A3 _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4730_ _1815_ _2157_ _2159_ immu_0.page_table\[15\]\[7\] _2167_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_56_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4661_ _2126_ _0753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6400_ _0782_ clknet_leaf_106_core_clock immu_0.page_table\[15\]\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3612_ _1309_ net685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6870__CLK clknet_leaf_67_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4592_ _2084_ _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_1501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_874 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6331_ _0713_ clknet_leaf_76_core_clock immu_1.page_table\[15\]\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3543_ _1271_ net557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6262_ _0644_ clknet_leaf_85_core_clock immu_1.page_table\[4\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3474_ _0906_ _1212_ _0912_ _1213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5856__A1 _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5213_ _2462_ _0160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6193_ _0575_ clknet_leaf_0_core_clock immu_0.page_table\[11\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_1253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5144_ _2419_ _0134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3253__C _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_2028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5459__I1 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6250__CLK clknet_leaf_83_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5075_ _2328_ _2367_ _2369_ immu_0.page_table\[8\]\[8\] _2378_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4026_ immu_1.page_table\[4\]\[9\] immu_1.page_table\[5\]\[9\] immu_1.page_table\[6\]\[9\]
+ immu_1.page_table\[7\]\[9\] _1441_ _1442_ _1687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__4831__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input202_I c1_sr_bus_data_o[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6033__A1 _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_2102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ net200 _2889_ _2891_ net956 _2905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4595__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3398__A2 _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4928_ net406 _2288_ _2289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_1989 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input98_I c0_sr_bus_data_o[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3709__B _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4859_ _2245_ _0023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4347__A1 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _0102_ clknet_leaf_8_core_clock immu_0.page_table\[8\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_12_core_clock_I clknet_3_3_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1077 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_2076 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_8_Left_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3173__I2 dmmu1.page_table\[14\]\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A2 _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6743__CLK clknet_leaf_39_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_2112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_944 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3228__I3 dmmu0.page_table\[7\]\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_1791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__B1 _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1887 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5838__A1 _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6273__CLK clknet_leaf_88_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3190_ _0936_ _0937_ _0938_ _0939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_0_79_1040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_2045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5900_ _2862_ _0447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6880_ _0453_ clknet_leaf_60_core_clock dmmu1.page_table\[7\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6015__A1 _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1011 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5831_ _2822_ _0418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4577__A1 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5762_ _2779_ _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_72_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1921 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4713_ _2156_ _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5693_ _2739_ _0363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4329__A1 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4204__I _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4644_ _2065_ _2108_ _2110_ net967 _2116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3248__C _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_2021 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_2032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4575_ _1838_ _1909_ _2028_ _2074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_12_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6616__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3526_ _1262_ net543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6314_ _0696_ clknet_leaf_96_core_clock dmmu1.page_table\[14\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_888 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_core_clock_I clknet_3_0_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6245_ _0627_ clknet_leaf_94_core_clock immu_1.page_table\[2\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3457_ _0896_ _1196_ _1197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input152_I c1_o_mem_high_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4501__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6176_ _3019_ _0566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6766__CLK clknet_leaf_31_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3388_ dmmu1.page_table\[4\]\[8\] dmmu1.page_table\[5\]\[8\] dmmu1.page_table\[6\]\[8\]
+ dmmu1.page_table\[7\]\[8\] _0898_ _0909_ _1130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_77_1725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5127_ _2408_ _0128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_78_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Right_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_1146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3068__A1 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5058_ _2368_ _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_58_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_1119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4265__B1 _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input13_I c0_o_mem_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4804__A2 _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_2036 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4009_ immu_0.page_table\[0\]\[8\] immu_0.page_table\[1\]\[8\] immu_0.page_table\[2\]\[8\]
+ immu_0.page_table\[3\]\[8\] _1487_ _1455_ _1671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_79_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4280__A3 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1032 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_871 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3091__I1 net23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_882 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4114__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5517__B1 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3791__A2 _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6296__CLK clknet_leaf_81_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_2394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3926__S0 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput310 ic0_wb_adr[10] net310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput321 ic0_wb_adr[6] net321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3846__A3 _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput332 ic1_mem_data[10] net332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput343 ic1_mem_data[20] net343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_1768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput354 ic1_mem_data[30] net354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7160__I net174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold50 dmmu0.page_table\[12\]\[12\] net784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput365 ic1_wb_adr[11] net365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold61 dmmu0.page_table\[11\]\[0\] net795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput376 ic1_wb_adr[7] net376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold72 dmmu0.page_table\[13\]\[11\] net806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput387 inner_wb_ack net387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold83 immu_1.page_table\[8\]\[1\] net817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput398 inner_wb_i_dat[3] net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3059__A1 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold94 immu_0.page_table\[9\]\[10\] net828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_3_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_2054 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_80_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3231__A1 _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6639__CLK clknet_leaf_25_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_917 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1949 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_3 net389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ _1940_ _0638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6789__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1083 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3311_ _0940_ _1055_ _0879_ _1056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_21_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4291_ _1851_ _1894_ _1897_ immu_1.page_table\[0\]\[3\] _1901_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5287__A2 _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6030_ _2935_ _0504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_56_1880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3242_ _0974_ _0979_ _0984_ _0988_ net523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_TAPCELL_ROW_56_1891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I c0_o_instr_long_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4495__B1 _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3173_ dmmu1.page_table\[12\]\[1\] dmmu1.page_table\[13\]\[1\] dmmu1.page_table\[14\]\[1\]
+ dmmu1.page_table\[15\]\[1\] _0908_ _0902_ _0922_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5039__A2 _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4798__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6932_ _0505_ clknet_leaf_58_core_clock dmmu1.page_table\[3\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3103__I _0854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5995__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6863_ _0436_ clknet_leaf_48_core_clock dmmu1.page_table\[8\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3470__A1 _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_2091 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_2053 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5814_ _2794_ _2802_ _2804_ net873 _2812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6794_ _0367_ clknet_leaf_49_core_clock dmmu1.page_table\[12\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_947 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3222__A1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5745_ _2769_ _0385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_50_1997 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_906 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5676_ _2059_ _2726_ _2728_ dmmu1.page_table\[13\]\[2\] _2731_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4627_ net198 _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3773__I _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4722__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input367_I ic1_wb_adr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4558_ _2063_ _2053_ _2055_ net943 _2064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_1161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3509_ net156 dmmu1.long_off_reg\[6\] _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4489_ _1852_ _2014_ _2016_ immu_1.page_table\[3\]\[3\] _2020_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_1178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _0610_ clknet_leaf_81_core_clock immu_1.page_table\[0\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3722__B _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6159_ _1863_ _3000_ _3002_ net945 _3010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_1539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1938 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5450__A2 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3300__I2 dmmu1.page_table\[14\]\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_869 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3461__A1 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5738__B1 _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output586_I net586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3213__A1 _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6931__CLK clknet_leaf_57_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6163__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7155__I net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_2445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_961 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_75_2467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1999 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5269__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput140 c1_o_mem_data[15] net140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput151 c1_o_mem_high_addr[1] net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput162 c1_o_mem_we net162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput173 c1_o_req_addr[3] net173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6311__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput184 c1_sr_bus_addr[12] net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput195 c1_sr_bus_addr[8] net195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4229__B1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_2031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_1038 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1937 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6461__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3860_ immu_0.page_table\[4\]\[4\] immu_0.page_table\[5\]\[4\] immu_0.page_table\[6\]\[4\]
+ immu_0.page_table\[7\]\[4\] _1396_ _1371_ _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_6_1183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3791_ _1382_ _1458_ _1375_ _1459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__4401__B1 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4952__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5530_ _2646_ _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_5_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5461_ immu_1.high_addr_off\[4\] _1855_ _2603_ _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7065__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4412_ _1970_ _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput603 net603 ic0_wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_23_972 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4704__A1 _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput614 net614 ic0_wb_i_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5392_ _1994_ _2552_ _2554_ dmmu0.page_table\[11\]\[11\] _2567_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_58_1942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5901__B1 _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput625 net625 ic1_mem_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput636 net636 ic1_mem_cache_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_2_877 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput647 net647 ic1_wb_i_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4343_ _1849_ _1927_ _1929_ net933 _1932_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7131_ net61 net584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_54_1817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput658 net658 inner_wb_4_burst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4180__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput669 net669 inner_wb_adr[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7062_ net300 net451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_10_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4274_ _1888_ _0604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_35_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6013_ _2776_ _2924_ _2926_ dmmu1.page_table\[3\]\[0\] _2927_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3225_ dmmu0.page_table\[12\]\[3\] dmmu0.page_table\[13\]\[3\] dmmu0.page_table\[14\]\[3\]
+ dmmu0.page_table\[15\]\[3\] _0950_ _0952_ _0972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_20_1075 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5680__A2 _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3156_ _0905_ _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_1717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_1859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3087_ net126 net21 _0842_ _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6804__CLK clknet_leaf_40_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input115_I c1_o_instr_long_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5432__A2 _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6915_ _0488_ clknet_leaf_54_core_clock dmmu1.page_table\[4\]\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4640__B1 _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1993 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6846_ _0419_ clknet_leaf_41_core_clock dmmu0.page_table\[1\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_1857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6954__CLK clknet_leaf_55_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6777_ _0350_ clknet_leaf_100_core_clock dmmu0.long_off_reg\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3989_ _1616_ _1649_ _1650_ _1651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_21_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5728_ _1826_ _1874_ _2031_ _2759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA_input80_I c0_sr_bus_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6145__B1 _3002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5659_ _2720_ _0348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold350 dmmu0.page_table\[12\]\[7\] net1084 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_70_2320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6334__CLK clknet_leaf_61_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4459__B1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5120__A1 _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_2064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_5_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1904 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output501_I net501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6484__CLK clknet_leaf_13_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5959__B1 _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_2135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2002 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_2046 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3985__A2 net241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_2079 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4934__A1 net407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_872 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_2518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_core_clock clknet_3_2_0_core_clock clknet_leaf_15_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_39_Left_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__B1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1031 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1064 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__CLK clknet_leaf_43_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4870__B1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6977__CLK clknet_leaf_103_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_1621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4961_ _2311_ _0059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3425__A1 _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4622__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6700_ _0273_ clknet_leaf_35_core_clock dmmu0.page_table\[4\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3912_ _1552_ _1576_ _1577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_28_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4892_ _1796_ _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_59_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_54_core_clock clknet_3_7_0_core_clock clknet_leaf_54_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_15_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5178__A1 _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6631_ _0204_ clknet_leaf_35_core_clock dmmu0.page_table\[12\]\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3843_ _1433_ _1506_ _1509_ _1434_ _1510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_6_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6207__CLK clknet_leaf_73_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3774_ immu_1.page_table\[4\]\[1\] immu_1.page_table\[5\]\[1\] immu_1.page_table\[6\]\[1\]
+ immu_1.page_table\[7\]\[1\] _1441_ _1442_ _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_27_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6562_ _0135_ clknet_leaf_20_core_clock immu_0.page_table\[5\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5513_ _2459_ _2630_ _2632_ dmmu0.page_table\[13\]\[5\] _2638_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6493_ _0066_ clknet_leaf_27_core_clock dmmu0.page_table\[14\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4212__I _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5444_ _1996_ _2581_ _2583_ net979 _2597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput411 net411 c0_i_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6357__CLK clknet_leaf_76_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput422 net422 c0_i_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput433 net433 c0_i_req_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_1240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5350__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput444 net444 c0_i_req_data[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4153__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput455 net455 c0_i_req_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5375_ _2558_ _0226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput466 net466 c1_i_mem_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7114_ net390 net567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput477 net477 c1_i_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput488 net488 c1_i_req_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4326_ _1921_ _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput499 net499 c1_i_req_data[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_17_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4257_ _1846_ _1876_ _1878_ net1051 _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7045_ net281 net432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input232_I dcache_wb_adr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3208_ dmmu0.page_table\[8\]\[2\] dmmu0.page_table\[9\]\[2\] dmmu0.page_table\[10\]\[2\]
+ dmmu0.page_table\[11\]\[2\] _0950_ _0952_ _0956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_78_1661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_1612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4188_ net197 _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_93_core_clock clknet_3_4_0_core_clock clknet_leaf_93_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3139_ _0888_ _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_1569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_942 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4613__B1 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1976 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_13_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6829_ _0402_ clknet_leaf_68_core_clock dmmu1.page_table\[10\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_2030 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6133__A3 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_2063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output451_I net451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1974 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold180 dmmu1.page_table\[6\]\[1\] net914 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold191 dmmu1.page_table\[3\]\[8\] net925 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5644__A2 _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3910__B _1574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1008 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3502__S1 net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4080__A1 _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_25_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__B1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1063 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4383__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_1858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3490_ _1180_ _1183_ _1228_ _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_64_1749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1017 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5332__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_36_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5160_ _2427_ _0142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_8_core_clock_I clknet_3_1_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4111_ icache_arbiter.o_sel_sig net379 _1766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5091_ _2269_ _2382_ _2384_ immu_0.page_table\[7\]\[3\] _2388_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_40_1760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4042_ immu_0.page_table\[4\]\[9\] immu_0.page_table\[5\]\[9\] immu_0.page_table\[6\]\[9\]
+ immu_0.page_table\[7\]\[9\] _1396_ _1371_ _1703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_79_1970 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3646__A1 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4843__B1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3741__S1 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1889 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5993_ _2790_ _2907_ _2909_ net1078 _2915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4944_ _2258_ _2299_ _2302_ dmmu0.page_table\[7\]\[0\] _2303_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_23_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4875_ _2253_ _0031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_1616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6614_ _0187_ clknet_leaf_5_core_clock immu_0.page_table\[0\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3826_ _1385_ immu_0.page_table\[14\]\[3\] _1493_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6545_ _0118_ clknet_leaf_18_core_clock immu_0.page_table\[7\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5571__A1 _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3757_ _1423_ _1425_ _1366_ _1426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input182_I c1_sr_bus_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _0049_ clknet_leaf_102_core_clock net406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_3688_ _1304_ _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4126__A2 _0815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5427_ _2588_ _0248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_1540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5874__A2 _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4098__B _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5358_ _2529_ _2536_ _2538_ net973 _2548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input43_I c0_o_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4309_ _1910_ _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5087__B1 _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5289_ _1805_ _2502_ _2504_ immu_0.page_table\[0\]\[4\] _2508_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5626__A2 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3637__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_2067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_1486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4062__A1 _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2005 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6522__CLK clknet_leaf_0_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4601__A3 _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_1451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output499_I net499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1940 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5011__B1 _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1984 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4365__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output666_I net666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_85_core_clock_I clknet_3_5_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6672__CLK clknet_leaf_33_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7163__I net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1891 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_1782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3420__S0 _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_2052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_1537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3100__I0 net132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5396__A4 _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_1259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_5_core_clock clknet_3_0_0_core_clock clknet_leaf_5_core_clock vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3800__A1 _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4660_ _2051_ _2123_ _2125_ immu_1.page_table\[11\]\[0\] _2126_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3239__S0 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3611_ _1308_ net256 _1309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5553__A1 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ _2067_ _2075_ _2077_ net1061 _2084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_40_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_981 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6330_ _0712_ clknet_leaf_71_core_clock immu_1.page_table\[15\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3542_ net148 net43 _1267_ _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1081 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5305__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6261_ _0643_ clknet_leaf_83_core_clock immu_1.page_table\[4\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_920 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_867 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3473_ dmmu1.page_table\[0\]\[11\] dmmu1.page_table\[1\]\[11\] dmmu1.page_table\[2\]\[11\]
+ dmmu1.page_table\[3\]\[11\] _0898_ _0901_ _1212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_10_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7073__I net357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_101_core_clock clknet_3_1_0_core_clock clknet_leaf_101_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_1991 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5856__A2 _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5212_ _2461_ _2447_ _2449_ immu_0.page_table\[3\]\[6\] _2462_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3867__A1 net5 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6192_ _0574_ clknet_leaf_1_core_clock immu_0.page_table\[11\]\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5143_ _2267_ _2414_ _2416_ net951 _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5069__B1 _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5608__A2 _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5074_ _2377_ _0106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3619__A1 _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4816__B1 _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4025_ immu_1.page_table\[0\]\[9\] immu_1.page_table\[1\]\[9\] immu_1.page_table\[2\]\[9\]
+ immu_1.page_table\[3\]\[9\] _1441_ _1442_ _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6545__CLK clknet_leaf_18_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6033__A2 _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5976_ _2904_ _0481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1962 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4927_ _1776_ _2285_ _2287_ _1823_ _2288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4595__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5792__A1 _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input397_I inner_wb_i_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4858_ _1777_ _2242_ _2244_ dmmu0.page_table\[9\]\[0\] _2245_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_1468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4347__A2 _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3809_ immu_1.page_table\[12\]\[2\] immu_1.page_table\[13\]\[2\] _1474_ _1477_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4789_ _2202_ _0805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_1722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6528_ _0101_ clknet_leaf_0_core_clock immu_0.page_table\[8\]\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_1154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3725__B _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1045 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_2071 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6459_ _0032_ clknet_leaf_12_core_clock dmmu0.page_table\[9\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1056 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1911 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1922 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_2088 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4283__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_901 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_912 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4035__A1 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1049 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5232__B1 _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_967 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7158__I net172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__A1 _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1866 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6418__CLK clknet_leaf_104_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5299__B1 _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4310__I _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5838__A2 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1052 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6568__CLK clknet_leaf_4_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1074 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_2040 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1085 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1902 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1913 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_2095 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_2057 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6015__A2 _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6173__S _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5830_ _1776_ _2819_ _2821_ net1019 _2822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_1258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5761_ _2682_ _2777_ _2779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7068__I net407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1067 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ _1790_ _2155_ _2156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_16_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5692_ _2105_ _2725_ _2727_ dmmu1.page_table\[13\]\[10\] _2739_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_907 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4329__A2 _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4643_ _2115_ _0746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4574_ _2073_ _0719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6313_ _0695_ clknet_leaf_94_core_clock immu_1.page_table\[3\]\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3525_ net134 net29 _0850_ _1262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_1327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4220__I _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6244_ _0626_ clknet_leaf_80_core_clock immu_1.page_table\[2\]\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3264__C _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3456_ dmmu1.page_table\[12\]\[10\] dmmu1.page_table\[13\]\[10\] dmmu1.page_table\[14\]\[10\]
+ dmmu1.page_table\[15\]\[10\] _0887_ _0900_ _1196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4501__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6175_ dmmu1.long_off_reg\[2\] _1849_ _3016_ _3019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3387_ dmmu1.page_table\[0\]\[8\] dmmu1.page_table\[1\]\[8\] dmmu1.page_table\[2\]\[8\]
+ dmmu1.page_table\[3\]\[8\] _0898_ _0909_ _1129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_1685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3560__I0 net161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input145_I c1_o_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5126_ _2277_ _2398_ _2400_ immu_0.page_table\[6\]\[7\] _2408_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_1950 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5057_ _2140_ _2366_ _2368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_2004 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4265__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3068__A2 _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input312_I ic0_wb_adr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4008_ immu_0.page_table\[4\]\[8\] immu_0.page_table\[5\]\[8\] immu_0.page_table\[6\]\[8\]
+ immu_0.page_table\[7\]\[8\] _1424_ _1455_ _1670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_75_1472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4017__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5959_ _2786_ _2890_ _2892_ net1074 _2896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_1191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3439__C _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5517__A1 _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1099 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_2384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6710__CLK clknet_leaf_26_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_2395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output629_I net629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput300 ic0_mem_data[30] net300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3926__S1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput311 ic0_wb_adr[11] net311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput322 ic0_wb_adr[7] net322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_1184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput333 ic1_mem_data[11] net333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput344 ic1_mem_data[21] net344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold40 immu_0.page_table\[4\]\[2\] net774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput355 ic1_mem_data[31] net355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold51 immu_0.page_table\[9\]\[7\] net785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold62 dmmu1.page_table\[12\]\[9\] net796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput366 ic1_wb_adr[12] net366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_26_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput377 ic1_wb_adr[8] net377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold73 immu_0.page_table\[6\]\[5\] net807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput388 inner_wb_err net388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput399 inner_wb_i_dat[4] net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3059__A2 _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold84 immu_0.page_table\[9\]\[9\] net818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6860__CLK clknet_leaf_47_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold95 dmmu0.page_table\[2\]\[1\] net829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_3_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1870 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1881 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5756__A1 _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1892 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3349__C _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3231__A2 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3862__S0 _1463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6240__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_20_Left_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_4 net389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1051 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5136__I _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3790__I0 _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3310_ dmmu0.page_table\[8\]\[5\] dmmu0.page_table\[9\]\[5\] dmmu0.page_table\[10\]\[5\]
+ dmmu0.page_table\[11\]\[5\] _0865_ _0868_ _1055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_10_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4290_ _1900_ _0608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6390__CLK clknet_leaf_80_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3241_ _0895_ _0987_ _0915_ _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_24_2094 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A1 _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3542__I0 net148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3172_ _0881_ _0885_ _0921_ _0822_ net520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_20_1235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5444__B1 _2583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6931_ _0504_ clknet_leaf_57_core_clock dmmu1.page_table\[3\]\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5995__A1 _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _0435_ clknet_leaf_48_core_clock dmmu1.page_table\[8\]\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1910 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5813_ _2811_ _0411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6793_ _0366_ clknet_leaf_45_core_clock dmmu1.page_table\[12\]\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1943 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5744_ _2067_ _2760_ _2762_ dmmu1.page_table\[11\]\[6\] _2769_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3853__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5675_ _2730_ _0354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_992 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4626_ _2104_ _0740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6733__CLK clknet_leaf_45_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4722__A2 _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_973 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4557_ _1854_ _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_input262_I dcache_wb_o_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3508_ _1119_ _1236_ _1245_ _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4488_ _2019_ _0687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6227_ _0609_ clknet_leaf_87_core_clock immu_1.page_table\[0\]\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3439_ _0878_ _1173_ _1178_ _0862_ _1179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4030__S0 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6883__CLK clknet_leaf_66_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3533__I0 net144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6158_ _3009_ _0558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5109_ _2397_ _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_38_1507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6089_ _2847_ _2958_ _2960_ net1082 _2969_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_68_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_11_Left_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3230__S _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3461__A2 _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5738__A1 _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_2063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6263__CLK clknet_leaf_86_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_2074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_24_core_clock_I clknet_3_2_0_core_clock vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_2571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_2582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6163__A1 _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_2457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1945 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1978 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3119__I3 dmmu0.page_table\[7\]\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7171__I net170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__A1 net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5674__B1 _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput130 c1_o_mem_addr[6] net130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput141 c1_o_mem_data[1] net141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput152 c1_o_mem_high_addr[2] net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_1022 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput163 c1_o_req_active net163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput174 c1_o_req_addr[4] net174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4229__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3204__I _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1044 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput185 c1_sr_bus_addr[13] net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5426__B1 _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput196 c1_sr_bus_addr[9] net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_1066 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1028 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5977__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6606__CLK clknet_leaf_15_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_2087 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1927 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_2098 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_1364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_44_core_clock clknet_3_6_0_core_clock clknet_leaf_44_core_clock vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_1651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_45_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4401__A1 _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3790_ _1456_ _1457_ _1377_ _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6756__CLK clknet_leaf_11_core_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_918 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4952__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_1747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5460_ _2607_ _0262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4411_ _1870_ _1956_ _1958_ immu_1.page_table\[6\]\[10\] _1970_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4165__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput604 net604 ic0_wb_i_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4704__A2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5901__A1 _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _2566_ _0234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput615 net615 ic0_wb_i_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_58_1943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput626 net626 ic1_mem_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7130_ net60 net583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput637 net637 ic1_mem_ppl_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_61_2069 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput648 net648 ic1_wb_i_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4342_ _1931_ _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput659 net659 inner_wb_8_burst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_39_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3823__B _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7061_ net298 net449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4273_ _1868_ _1876_ _1878_ immu_1.page_table\[7\]\[9\] _1888_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6012_ _2925_ _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3224_ dmmu0.page_table\[8\]\[3\] dmmu0.page_table\[9\]\[3\] dmmu0.page_table\[10\]\[3\]
+ dmmu0.page_table\[11\]\[3\] _0950_ _0948_ _0971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
.ends

