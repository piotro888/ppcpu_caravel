magic
tech sky130A
magscale 1 2
timestamp 1672421699
<< obsli1 >>
rect 1104 2159 58880 157777
<< obsm1 >>
rect 566 1912 59970 157808
<< metal2 >>
rect 1398 0 1454 800
rect 2226 0 2282 800
rect 3054 0 3110 800
rect 3882 0 3938 800
rect 4710 0 4766 800
rect 5538 0 5594 800
rect 6366 0 6422 800
rect 7194 0 7250 800
rect 8022 0 8078 800
rect 8850 0 8906 800
rect 9678 0 9734 800
rect 10506 0 10562 800
rect 11334 0 11390 800
rect 12162 0 12218 800
rect 12990 0 13046 800
rect 13818 0 13874 800
rect 14646 0 14702 800
rect 15474 0 15530 800
rect 16302 0 16358 800
rect 17130 0 17186 800
rect 17958 0 18014 800
rect 18786 0 18842 800
rect 19614 0 19670 800
rect 20442 0 20498 800
rect 21270 0 21326 800
rect 22098 0 22154 800
rect 22926 0 22982 800
rect 23754 0 23810 800
rect 24582 0 24638 800
rect 25410 0 25466 800
rect 26238 0 26294 800
rect 27066 0 27122 800
rect 27894 0 27950 800
rect 28722 0 28778 800
rect 29550 0 29606 800
rect 30378 0 30434 800
rect 31206 0 31262 800
rect 32034 0 32090 800
rect 32862 0 32918 800
rect 33690 0 33746 800
rect 34518 0 34574 800
rect 35346 0 35402 800
rect 36174 0 36230 800
rect 37002 0 37058 800
rect 37830 0 37886 800
rect 38658 0 38714 800
rect 39486 0 39542 800
rect 40314 0 40370 800
rect 41142 0 41198 800
rect 41970 0 42026 800
rect 42798 0 42854 800
rect 43626 0 43682 800
rect 44454 0 44510 800
rect 45282 0 45338 800
rect 46110 0 46166 800
rect 46938 0 46994 800
rect 47766 0 47822 800
rect 48594 0 48650 800
rect 49422 0 49478 800
rect 50250 0 50306 800
rect 51078 0 51134 800
rect 51906 0 51962 800
rect 52734 0 52790 800
rect 53562 0 53618 800
rect 54390 0 54446 800
rect 55218 0 55274 800
rect 56046 0 56102 800
rect 56874 0 56930 800
rect 57702 0 57758 800
rect 58530 0 58586 800
<< obsm2 >>
rect 572 856 59964 157797
rect 572 800 1342 856
rect 1510 800 2170 856
rect 2338 800 2998 856
rect 3166 800 3826 856
rect 3994 800 4654 856
rect 4822 800 5482 856
rect 5650 800 6310 856
rect 6478 800 7138 856
rect 7306 800 7966 856
rect 8134 800 8794 856
rect 8962 800 9622 856
rect 9790 800 10450 856
rect 10618 800 11278 856
rect 11446 800 12106 856
rect 12274 800 12934 856
rect 13102 800 13762 856
rect 13930 800 14590 856
rect 14758 800 15418 856
rect 15586 800 16246 856
rect 16414 800 17074 856
rect 17242 800 17902 856
rect 18070 800 18730 856
rect 18898 800 19558 856
rect 19726 800 20386 856
rect 20554 800 21214 856
rect 21382 800 22042 856
rect 22210 800 22870 856
rect 23038 800 23698 856
rect 23866 800 24526 856
rect 24694 800 25354 856
rect 25522 800 26182 856
rect 26350 800 27010 856
rect 27178 800 27838 856
rect 28006 800 28666 856
rect 28834 800 29494 856
rect 29662 800 30322 856
rect 30490 800 31150 856
rect 31318 800 31978 856
rect 32146 800 32806 856
rect 32974 800 33634 856
rect 33802 800 34462 856
rect 34630 800 35290 856
rect 35458 800 36118 856
rect 36286 800 36946 856
rect 37114 800 37774 856
rect 37942 800 38602 856
rect 38770 800 39430 856
rect 39598 800 40258 856
rect 40426 800 41086 856
rect 41254 800 41914 856
rect 42082 800 42742 856
rect 42910 800 43570 856
rect 43738 800 44398 856
rect 44566 800 45226 856
rect 45394 800 46054 856
rect 46222 800 46882 856
rect 47050 800 47710 856
rect 47878 800 48538 856
rect 48706 800 49366 856
rect 49534 800 50194 856
rect 50362 800 51022 856
rect 51190 800 51850 856
rect 52018 800 52678 856
rect 52846 800 53506 856
rect 53674 800 54334 856
rect 54502 800 55162 856
rect 55330 800 55990 856
rect 56158 800 56818 856
rect 56986 800 57646 856
rect 57814 800 58474 856
rect 58642 800 59964 856
<< metal3 >>
rect 59200 143896 60000 144016
rect 59200 143488 60000 143608
rect 59200 143080 60000 143200
rect 59200 142672 60000 142792
rect 59200 142264 60000 142384
rect 59200 141856 60000 141976
rect 59200 141448 60000 141568
rect 59200 141040 60000 141160
rect 59200 140632 60000 140752
rect 59200 140224 60000 140344
rect 59200 139816 60000 139936
rect 59200 139408 60000 139528
rect 59200 139000 60000 139120
rect 59200 138592 60000 138712
rect 59200 138184 60000 138304
rect 59200 137776 60000 137896
rect 0 137368 800 137488
rect 59200 137368 60000 137488
rect 0 137096 800 137216
rect 0 136824 800 136944
rect 59200 136960 60000 137080
rect 0 136552 800 136672
rect 59200 136552 60000 136672
rect 0 136280 800 136400
rect 0 136008 800 136128
rect 59200 136144 60000 136264
rect 0 135736 800 135856
rect 59200 135736 60000 135856
rect 0 135464 800 135584
rect 0 135192 800 135312
rect 59200 135328 60000 135448
rect 0 134920 800 135040
rect 59200 134920 60000 135040
rect 0 134648 800 134768
rect 0 134376 800 134496
rect 59200 134512 60000 134632
rect 0 134104 800 134224
rect 59200 134104 60000 134224
rect 0 133832 800 133952
rect 0 133560 800 133680
rect 59200 133696 60000 133816
rect 0 133288 800 133408
rect 59200 133288 60000 133408
rect 0 133016 800 133136
rect 0 132744 800 132864
rect 59200 132880 60000 133000
rect 0 132472 800 132592
rect 59200 132472 60000 132592
rect 0 132200 800 132320
rect 0 131928 800 132048
rect 59200 132064 60000 132184
rect 0 131656 800 131776
rect 59200 131656 60000 131776
rect 0 131384 800 131504
rect 0 131112 800 131232
rect 59200 131248 60000 131368
rect 0 130840 800 130960
rect 59200 130840 60000 130960
rect 0 130568 800 130688
rect 0 130296 800 130416
rect 59200 130432 60000 130552
rect 0 130024 800 130144
rect 59200 130024 60000 130144
rect 0 129752 800 129872
rect 0 129480 800 129600
rect 59200 129616 60000 129736
rect 0 129208 800 129328
rect 59200 129208 60000 129328
rect 0 128936 800 129056
rect 0 128664 800 128784
rect 59200 128800 60000 128920
rect 0 128392 800 128512
rect 59200 128392 60000 128512
rect 0 128120 800 128240
rect 0 127848 800 127968
rect 59200 127984 60000 128104
rect 0 127576 800 127696
rect 59200 127576 60000 127696
rect 0 127304 800 127424
rect 0 127032 800 127152
rect 59200 127168 60000 127288
rect 0 126760 800 126880
rect 59200 126760 60000 126880
rect 0 126488 800 126608
rect 0 126216 800 126336
rect 59200 126352 60000 126472
rect 0 125944 800 126064
rect 59200 125944 60000 126064
rect 0 125672 800 125792
rect 0 125400 800 125520
rect 59200 125536 60000 125656
rect 0 125128 800 125248
rect 59200 125128 60000 125248
rect 0 124856 800 124976
rect 0 124584 800 124704
rect 59200 124720 60000 124840
rect 0 124312 800 124432
rect 59200 124312 60000 124432
rect 0 124040 800 124160
rect 0 123768 800 123888
rect 59200 123904 60000 124024
rect 0 123496 800 123616
rect 59200 123496 60000 123616
rect 0 123224 800 123344
rect 0 122952 800 123072
rect 59200 123088 60000 123208
rect 0 122680 800 122800
rect 59200 122680 60000 122800
rect 0 122408 800 122528
rect 0 122136 800 122256
rect 59200 122272 60000 122392
rect 0 121864 800 121984
rect 59200 121864 60000 121984
rect 0 121592 800 121712
rect 0 121320 800 121440
rect 59200 121456 60000 121576
rect 0 121048 800 121168
rect 59200 121048 60000 121168
rect 0 120776 800 120896
rect 0 120504 800 120624
rect 59200 120640 60000 120760
rect 0 120232 800 120352
rect 59200 120232 60000 120352
rect 0 119960 800 120080
rect 0 119688 800 119808
rect 59200 119824 60000 119944
rect 0 119416 800 119536
rect 59200 119416 60000 119536
rect 0 119144 800 119264
rect 0 118872 800 118992
rect 59200 119008 60000 119128
rect 0 118600 800 118720
rect 59200 118600 60000 118720
rect 0 118328 800 118448
rect 0 118056 800 118176
rect 59200 118192 60000 118312
rect 0 117784 800 117904
rect 59200 117784 60000 117904
rect 0 117512 800 117632
rect 0 117240 800 117360
rect 59200 117376 60000 117496
rect 0 116968 800 117088
rect 59200 116968 60000 117088
rect 0 116696 800 116816
rect 0 116424 800 116544
rect 59200 116560 60000 116680
rect 0 116152 800 116272
rect 59200 116152 60000 116272
rect 0 115880 800 116000
rect 0 115608 800 115728
rect 59200 115744 60000 115864
rect 0 115336 800 115456
rect 59200 115336 60000 115456
rect 0 115064 800 115184
rect 0 114792 800 114912
rect 59200 114928 60000 115048
rect 0 114520 800 114640
rect 59200 114520 60000 114640
rect 0 114248 800 114368
rect 0 113976 800 114096
rect 59200 114112 60000 114232
rect 0 113704 800 113824
rect 59200 113704 60000 113824
rect 0 113432 800 113552
rect 0 113160 800 113280
rect 59200 113296 60000 113416
rect 0 112888 800 113008
rect 59200 112888 60000 113008
rect 0 112616 800 112736
rect 0 112344 800 112464
rect 59200 112480 60000 112600
rect 0 112072 800 112192
rect 59200 112072 60000 112192
rect 0 111800 800 111920
rect 0 111528 800 111648
rect 59200 111664 60000 111784
rect 0 111256 800 111376
rect 59200 111256 60000 111376
rect 0 110984 800 111104
rect 0 110712 800 110832
rect 59200 110848 60000 110968
rect 0 110440 800 110560
rect 59200 110440 60000 110560
rect 0 110168 800 110288
rect 0 109896 800 110016
rect 59200 110032 60000 110152
rect 0 109624 800 109744
rect 59200 109624 60000 109744
rect 0 109352 800 109472
rect 0 109080 800 109200
rect 59200 109216 60000 109336
rect 0 108808 800 108928
rect 59200 108808 60000 108928
rect 0 108536 800 108656
rect 0 108264 800 108384
rect 59200 108400 60000 108520
rect 0 107992 800 108112
rect 59200 107992 60000 108112
rect 0 107720 800 107840
rect 0 107448 800 107568
rect 59200 107584 60000 107704
rect 0 107176 800 107296
rect 59200 107176 60000 107296
rect 0 106904 800 107024
rect 0 106632 800 106752
rect 59200 106768 60000 106888
rect 0 106360 800 106480
rect 59200 106360 60000 106480
rect 0 106088 800 106208
rect 0 105816 800 105936
rect 59200 105952 60000 106072
rect 0 105544 800 105664
rect 59200 105544 60000 105664
rect 0 105272 800 105392
rect 0 105000 800 105120
rect 59200 105136 60000 105256
rect 0 104728 800 104848
rect 59200 104728 60000 104848
rect 0 104456 800 104576
rect 0 104184 800 104304
rect 59200 104320 60000 104440
rect 0 103912 800 104032
rect 59200 103912 60000 104032
rect 0 103640 800 103760
rect 0 103368 800 103488
rect 59200 103504 60000 103624
rect 0 103096 800 103216
rect 59200 103096 60000 103216
rect 0 102824 800 102944
rect 0 102552 800 102672
rect 59200 102688 60000 102808
rect 0 102280 800 102400
rect 59200 102280 60000 102400
rect 0 102008 800 102128
rect 0 101736 800 101856
rect 59200 101872 60000 101992
rect 0 101464 800 101584
rect 59200 101464 60000 101584
rect 0 101192 800 101312
rect 0 100920 800 101040
rect 59200 101056 60000 101176
rect 0 100648 800 100768
rect 59200 100648 60000 100768
rect 0 100376 800 100496
rect 0 100104 800 100224
rect 59200 100240 60000 100360
rect 0 99832 800 99952
rect 59200 99832 60000 99952
rect 0 99560 800 99680
rect 0 99288 800 99408
rect 59200 99424 60000 99544
rect 0 99016 800 99136
rect 59200 99016 60000 99136
rect 0 98744 800 98864
rect 0 98472 800 98592
rect 59200 98608 60000 98728
rect 0 98200 800 98320
rect 59200 98200 60000 98320
rect 0 97928 800 98048
rect 0 97656 800 97776
rect 59200 97792 60000 97912
rect 0 97384 800 97504
rect 59200 97384 60000 97504
rect 0 97112 800 97232
rect 0 96840 800 96960
rect 59200 96976 60000 97096
rect 0 96568 800 96688
rect 59200 96568 60000 96688
rect 0 96296 800 96416
rect 0 96024 800 96144
rect 59200 96160 60000 96280
rect 0 95752 800 95872
rect 59200 95752 60000 95872
rect 0 95480 800 95600
rect 0 95208 800 95328
rect 59200 95344 60000 95464
rect 0 94936 800 95056
rect 59200 94936 60000 95056
rect 0 94664 800 94784
rect 0 94392 800 94512
rect 59200 94528 60000 94648
rect 0 94120 800 94240
rect 59200 94120 60000 94240
rect 0 93848 800 93968
rect 0 93576 800 93696
rect 59200 93712 60000 93832
rect 0 93304 800 93424
rect 59200 93304 60000 93424
rect 0 93032 800 93152
rect 0 92760 800 92880
rect 59200 92896 60000 93016
rect 0 92488 800 92608
rect 59200 92488 60000 92608
rect 0 92216 800 92336
rect 0 91944 800 92064
rect 59200 92080 60000 92200
rect 0 91672 800 91792
rect 59200 91672 60000 91792
rect 0 91400 800 91520
rect 0 91128 800 91248
rect 59200 91264 60000 91384
rect 0 90856 800 90976
rect 59200 90856 60000 90976
rect 0 90584 800 90704
rect 0 90312 800 90432
rect 59200 90448 60000 90568
rect 0 90040 800 90160
rect 59200 90040 60000 90160
rect 0 89768 800 89888
rect 0 89496 800 89616
rect 59200 89632 60000 89752
rect 0 89224 800 89344
rect 59200 89224 60000 89344
rect 0 88952 800 89072
rect 0 88680 800 88800
rect 59200 88816 60000 88936
rect 0 88408 800 88528
rect 59200 88408 60000 88528
rect 0 88136 800 88256
rect 0 87864 800 87984
rect 59200 88000 60000 88120
rect 0 87592 800 87712
rect 59200 87592 60000 87712
rect 0 87320 800 87440
rect 0 87048 800 87168
rect 59200 87184 60000 87304
rect 0 86776 800 86896
rect 59200 86776 60000 86896
rect 0 86504 800 86624
rect 0 86232 800 86352
rect 59200 86368 60000 86488
rect 0 85960 800 86080
rect 59200 85960 60000 86080
rect 0 85688 800 85808
rect 0 85416 800 85536
rect 59200 85552 60000 85672
rect 0 85144 800 85264
rect 59200 85144 60000 85264
rect 0 84872 800 84992
rect 0 84600 800 84720
rect 59200 84736 60000 84856
rect 0 84328 800 84448
rect 59200 84328 60000 84448
rect 0 84056 800 84176
rect 0 83784 800 83904
rect 59200 83920 60000 84040
rect 0 83512 800 83632
rect 59200 83512 60000 83632
rect 0 83240 800 83360
rect 0 82968 800 83088
rect 59200 83104 60000 83224
rect 0 82696 800 82816
rect 59200 82696 60000 82816
rect 0 82424 800 82544
rect 0 82152 800 82272
rect 59200 82288 60000 82408
rect 0 81880 800 82000
rect 59200 81880 60000 82000
rect 0 81608 800 81728
rect 0 81336 800 81456
rect 59200 81472 60000 81592
rect 0 81064 800 81184
rect 59200 81064 60000 81184
rect 0 80792 800 80912
rect 0 80520 800 80640
rect 59200 80656 60000 80776
rect 0 80248 800 80368
rect 59200 80248 60000 80368
rect 0 79976 800 80096
rect 0 79704 800 79824
rect 59200 79840 60000 79960
rect 0 79432 800 79552
rect 59200 79432 60000 79552
rect 0 79160 800 79280
rect 0 78888 800 79008
rect 59200 79024 60000 79144
rect 0 78616 800 78736
rect 59200 78616 60000 78736
rect 0 78344 800 78464
rect 0 78072 800 78192
rect 59200 78208 60000 78328
rect 0 77800 800 77920
rect 59200 77800 60000 77920
rect 0 77528 800 77648
rect 0 77256 800 77376
rect 59200 77392 60000 77512
rect 0 76984 800 77104
rect 59200 76984 60000 77104
rect 0 76712 800 76832
rect 0 76440 800 76560
rect 59200 76576 60000 76696
rect 0 76168 800 76288
rect 59200 76168 60000 76288
rect 0 75896 800 76016
rect 0 75624 800 75744
rect 59200 75760 60000 75880
rect 0 75352 800 75472
rect 59200 75352 60000 75472
rect 0 75080 800 75200
rect 0 74808 800 74928
rect 59200 74944 60000 75064
rect 0 74536 800 74656
rect 59200 74536 60000 74656
rect 0 74264 800 74384
rect 0 73992 800 74112
rect 59200 74128 60000 74248
rect 0 73720 800 73840
rect 59200 73720 60000 73840
rect 0 73448 800 73568
rect 0 73176 800 73296
rect 59200 73312 60000 73432
rect 0 72904 800 73024
rect 59200 72904 60000 73024
rect 0 72632 800 72752
rect 0 72360 800 72480
rect 59200 72496 60000 72616
rect 0 72088 800 72208
rect 59200 72088 60000 72208
rect 0 71816 800 71936
rect 0 71544 800 71664
rect 59200 71680 60000 71800
rect 0 71272 800 71392
rect 59200 71272 60000 71392
rect 0 71000 800 71120
rect 0 70728 800 70848
rect 59200 70864 60000 70984
rect 0 70456 800 70576
rect 59200 70456 60000 70576
rect 0 70184 800 70304
rect 0 69912 800 70032
rect 59200 70048 60000 70168
rect 0 69640 800 69760
rect 59200 69640 60000 69760
rect 0 69368 800 69488
rect 0 69096 800 69216
rect 59200 69232 60000 69352
rect 0 68824 800 68944
rect 59200 68824 60000 68944
rect 0 68552 800 68672
rect 0 68280 800 68400
rect 59200 68416 60000 68536
rect 0 68008 800 68128
rect 59200 68008 60000 68128
rect 0 67736 800 67856
rect 0 67464 800 67584
rect 59200 67600 60000 67720
rect 0 67192 800 67312
rect 59200 67192 60000 67312
rect 0 66920 800 67040
rect 0 66648 800 66768
rect 59200 66784 60000 66904
rect 0 66376 800 66496
rect 59200 66376 60000 66496
rect 0 66104 800 66224
rect 0 65832 800 65952
rect 59200 65968 60000 66088
rect 0 65560 800 65680
rect 59200 65560 60000 65680
rect 0 65288 800 65408
rect 0 65016 800 65136
rect 59200 65152 60000 65272
rect 0 64744 800 64864
rect 59200 64744 60000 64864
rect 0 64472 800 64592
rect 0 64200 800 64320
rect 59200 64336 60000 64456
rect 0 63928 800 64048
rect 59200 63928 60000 64048
rect 0 63656 800 63776
rect 0 63384 800 63504
rect 59200 63520 60000 63640
rect 0 63112 800 63232
rect 59200 63112 60000 63232
rect 0 62840 800 62960
rect 0 62568 800 62688
rect 59200 62704 60000 62824
rect 0 62296 800 62416
rect 59200 62296 60000 62416
rect 0 62024 800 62144
rect 0 61752 800 61872
rect 59200 61888 60000 62008
rect 0 61480 800 61600
rect 59200 61480 60000 61600
rect 0 61208 800 61328
rect 0 60936 800 61056
rect 59200 61072 60000 61192
rect 0 60664 800 60784
rect 59200 60664 60000 60784
rect 0 60392 800 60512
rect 0 60120 800 60240
rect 59200 60256 60000 60376
rect 0 59848 800 59968
rect 59200 59848 60000 59968
rect 0 59576 800 59696
rect 0 59304 800 59424
rect 59200 59440 60000 59560
rect 0 59032 800 59152
rect 59200 59032 60000 59152
rect 0 58760 800 58880
rect 0 58488 800 58608
rect 59200 58624 60000 58744
rect 0 58216 800 58336
rect 59200 58216 60000 58336
rect 0 57944 800 58064
rect 0 57672 800 57792
rect 59200 57808 60000 57928
rect 0 57400 800 57520
rect 59200 57400 60000 57520
rect 0 57128 800 57248
rect 0 56856 800 56976
rect 59200 56992 60000 57112
rect 0 56584 800 56704
rect 59200 56584 60000 56704
rect 0 56312 800 56432
rect 0 56040 800 56160
rect 59200 56176 60000 56296
rect 0 55768 800 55888
rect 59200 55768 60000 55888
rect 0 55496 800 55616
rect 0 55224 800 55344
rect 59200 55360 60000 55480
rect 0 54952 800 55072
rect 59200 54952 60000 55072
rect 0 54680 800 54800
rect 0 54408 800 54528
rect 59200 54544 60000 54664
rect 0 54136 800 54256
rect 59200 54136 60000 54256
rect 0 53864 800 53984
rect 0 53592 800 53712
rect 59200 53728 60000 53848
rect 0 53320 800 53440
rect 59200 53320 60000 53440
rect 0 53048 800 53168
rect 0 52776 800 52896
rect 59200 52912 60000 53032
rect 0 52504 800 52624
rect 59200 52504 60000 52624
rect 0 52232 800 52352
rect 0 51960 800 52080
rect 59200 52096 60000 52216
rect 0 51688 800 51808
rect 59200 51688 60000 51808
rect 0 51416 800 51536
rect 0 51144 800 51264
rect 59200 51280 60000 51400
rect 0 50872 800 50992
rect 59200 50872 60000 50992
rect 0 50600 800 50720
rect 0 50328 800 50448
rect 59200 50464 60000 50584
rect 0 50056 800 50176
rect 59200 50056 60000 50176
rect 0 49784 800 49904
rect 0 49512 800 49632
rect 59200 49648 60000 49768
rect 0 49240 800 49360
rect 59200 49240 60000 49360
rect 0 48968 800 49088
rect 0 48696 800 48816
rect 59200 48832 60000 48952
rect 0 48424 800 48544
rect 59200 48424 60000 48544
rect 0 48152 800 48272
rect 0 47880 800 48000
rect 59200 48016 60000 48136
rect 0 47608 800 47728
rect 59200 47608 60000 47728
rect 0 47336 800 47456
rect 0 47064 800 47184
rect 59200 47200 60000 47320
rect 0 46792 800 46912
rect 59200 46792 60000 46912
rect 0 46520 800 46640
rect 0 46248 800 46368
rect 59200 46384 60000 46504
rect 0 45976 800 46096
rect 59200 45976 60000 46096
rect 0 45704 800 45824
rect 0 45432 800 45552
rect 59200 45568 60000 45688
rect 0 45160 800 45280
rect 59200 45160 60000 45280
rect 0 44888 800 45008
rect 0 44616 800 44736
rect 59200 44752 60000 44872
rect 0 44344 800 44464
rect 59200 44344 60000 44464
rect 0 44072 800 44192
rect 0 43800 800 43920
rect 59200 43936 60000 44056
rect 0 43528 800 43648
rect 59200 43528 60000 43648
rect 0 43256 800 43376
rect 0 42984 800 43104
rect 59200 43120 60000 43240
rect 0 42712 800 42832
rect 59200 42712 60000 42832
rect 0 42440 800 42560
rect 0 42168 800 42288
rect 59200 42304 60000 42424
rect 0 41896 800 42016
rect 59200 41896 60000 42016
rect 0 41624 800 41744
rect 0 41352 800 41472
rect 59200 41488 60000 41608
rect 0 41080 800 41200
rect 59200 41080 60000 41200
rect 0 40808 800 40928
rect 0 40536 800 40656
rect 59200 40672 60000 40792
rect 0 40264 800 40384
rect 59200 40264 60000 40384
rect 0 39992 800 40112
rect 0 39720 800 39840
rect 59200 39856 60000 39976
rect 0 39448 800 39568
rect 59200 39448 60000 39568
rect 0 39176 800 39296
rect 0 38904 800 39024
rect 59200 39040 60000 39160
rect 0 38632 800 38752
rect 59200 38632 60000 38752
rect 0 38360 800 38480
rect 0 38088 800 38208
rect 59200 38224 60000 38344
rect 0 37816 800 37936
rect 59200 37816 60000 37936
rect 0 37544 800 37664
rect 0 37272 800 37392
rect 59200 37408 60000 37528
rect 0 37000 800 37120
rect 59200 37000 60000 37120
rect 0 36728 800 36848
rect 0 36456 800 36576
rect 59200 36592 60000 36712
rect 0 36184 800 36304
rect 59200 36184 60000 36304
rect 0 35912 800 36032
rect 0 35640 800 35760
rect 59200 35776 60000 35896
rect 0 35368 800 35488
rect 59200 35368 60000 35488
rect 0 35096 800 35216
rect 0 34824 800 34944
rect 59200 34960 60000 35080
rect 0 34552 800 34672
rect 59200 34552 60000 34672
rect 0 34280 800 34400
rect 0 34008 800 34128
rect 59200 34144 60000 34264
rect 0 33736 800 33856
rect 59200 33736 60000 33856
rect 0 33464 800 33584
rect 0 33192 800 33312
rect 59200 33328 60000 33448
rect 0 32920 800 33040
rect 59200 32920 60000 33040
rect 0 32648 800 32768
rect 0 32376 800 32496
rect 59200 32512 60000 32632
rect 0 32104 800 32224
rect 59200 32104 60000 32224
rect 0 31832 800 31952
rect 0 31560 800 31680
rect 59200 31696 60000 31816
rect 0 31288 800 31408
rect 59200 31288 60000 31408
rect 0 31016 800 31136
rect 0 30744 800 30864
rect 59200 30880 60000 31000
rect 0 30472 800 30592
rect 59200 30472 60000 30592
rect 0 30200 800 30320
rect 0 29928 800 30048
rect 59200 30064 60000 30184
rect 0 29656 800 29776
rect 59200 29656 60000 29776
rect 0 29384 800 29504
rect 0 29112 800 29232
rect 59200 29248 60000 29368
rect 0 28840 800 28960
rect 59200 28840 60000 28960
rect 0 28568 800 28688
rect 0 28296 800 28416
rect 59200 28432 60000 28552
rect 0 28024 800 28144
rect 59200 28024 60000 28144
rect 0 27752 800 27872
rect 0 27480 800 27600
rect 59200 27616 60000 27736
rect 0 27208 800 27328
rect 59200 27208 60000 27328
rect 0 26936 800 27056
rect 0 26664 800 26784
rect 59200 26800 60000 26920
rect 0 26392 800 26512
rect 59200 26392 60000 26512
rect 0 26120 800 26240
rect 0 25848 800 25968
rect 59200 25984 60000 26104
rect 0 25576 800 25696
rect 59200 25576 60000 25696
rect 0 25304 800 25424
rect 0 25032 800 25152
rect 59200 25168 60000 25288
rect 0 24760 800 24880
rect 59200 24760 60000 24880
rect 0 24488 800 24608
rect 0 24216 800 24336
rect 59200 24352 60000 24472
rect 0 23944 800 24064
rect 59200 23944 60000 24064
rect 0 23672 800 23792
rect 0 23400 800 23520
rect 59200 23536 60000 23656
rect 0 23128 800 23248
rect 59200 23128 60000 23248
rect 0 22856 800 22976
rect 0 22584 800 22704
rect 59200 22720 60000 22840
rect 0 22312 800 22432
rect 59200 22312 60000 22432
rect 59200 21904 60000 22024
rect 59200 21496 60000 21616
rect 59200 21088 60000 21208
rect 59200 20680 60000 20800
rect 59200 20272 60000 20392
rect 59200 19864 60000 19984
rect 59200 19456 60000 19576
rect 59200 19048 60000 19168
rect 59200 18640 60000 18760
rect 59200 18232 60000 18352
rect 59200 17824 60000 17944
rect 59200 17416 60000 17536
rect 59200 17008 60000 17128
rect 59200 16600 60000 16720
rect 59200 16192 60000 16312
rect 59200 15784 60000 15904
<< obsm3 >>
rect 800 144096 59200 157793
rect 800 143816 59120 144096
rect 800 143688 59200 143816
rect 800 143408 59120 143688
rect 800 143280 59200 143408
rect 800 143000 59120 143280
rect 800 142872 59200 143000
rect 800 142592 59120 142872
rect 800 142464 59200 142592
rect 800 142184 59120 142464
rect 800 142056 59200 142184
rect 800 141776 59120 142056
rect 800 141648 59200 141776
rect 800 141368 59120 141648
rect 800 141240 59200 141368
rect 800 140960 59120 141240
rect 800 140832 59200 140960
rect 800 140552 59120 140832
rect 800 140424 59200 140552
rect 800 140144 59120 140424
rect 800 140016 59200 140144
rect 800 139736 59120 140016
rect 800 139608 59200 139736
rect 800 139328 59120 139608
rect 800 139200 59200 139328
rect 800 138920 59120 139200
rect 800 138792 59200 138920
rect 800 138512 59120 138792
rect 800 138384 59200 138512
rect 800 138104 59120 138384
rect 800 137976 59200 138104
rect 800 137696 59120 137976
rect 800 137568 59200 137696
rect 880 137288 59120 137568
rect 880 137160 59200 137288
rect 880 136880 59120 137160
rect 880 136752 59200 136880
rect 880 136472 59120 136752
rect 880 136344 59200 136472
rect 880 136064 59120 136344
rect 880 135936 59200 136064
rect 880 135656 59120 135936
rect 880 135528 59200 135656
rect 880 135248 59120 135528
rect 880 135120 59200 135248
rect 880 134840 59120 135120
rect 880 134712 59200 134840
rect 880 134432 59120 134712
rect 880 134304 59200 134432
rect 880 134024 59120 134304
rect 880 133896 59200 134024
rect 880 133616 59120 133896
rect 880 133488 59200 133616
rect 880 133208 59120 133488
rect 880 133080 59200 133208
rect 880 132800 59120 133080
rect 880 132672 59200 132800
rect 880 132392 59120 132672
rect 880 132264 59200 132392
rect 880 131984 59120 132264
rect 880 131856 59200 131984
rect 880 131576 59120 131856
rect 880 131448 59200 131576
rect 880 131168 59120 131448
rect 880 131040 59200 131168
rect 880 130760 59120 131040
rect 880 130632 59200 130760
rect 880 130352 59120 130632
rect 880 130224 59200 130352
rect 880 129944 59120 130224
rect 880 129816 59200 129944
rect 880 129536 59120 129816
rect 880 129408 59200 129536
rect 880 129128 59120 129408
rect 880 129000 59200 129128
rect 880 128720 59120 129000
rect 880 128592 59200 128720
rect 880 128312 59120 128592
rect 880 128184 59200 128312
rect 880 127904 59120 128184
rect 880 127776 59200 127904
rect 880 127496 59120 127776
rect 880 127368 59200 127496
rect 880 127088 59120 127368
rect 880 126960 59200 127088
rect 880 126680 59120 126960
rect 880 126552 59200 126680
rect 880 126272 59120 126552
rect 880 126144 59200 126272
rect 880 125864 59120 126144
rect 880 125736 59200 125864
rect 880 125456 59120 125736
rect 880 125328 59200 125456
rect 880 125048 59120 125328
rect 880 124920 59200 125048
rect 880 124640 59120 124920
rect 880 124512 59200 124640
rect 880 124232 59120 124512
rect 880 124104 59200 124232
rect 880 123824 59120 124104
rect 880 123696 59200 123824
rect 880 123416 59120 123696
rect 880 123288 59200 123416
rect 880 123008 59120 123288
rect 880 122880 59200 123008
rect 880 122600 59120 122880
rect 880 122472 59200 122600
rect 880 122192 59120 122472
rect 880 122064 59200 122192
rect 880 121784 59120 122064
rect 880 121656 59200 121784
rect 880 121376 59120 121656
rect 880 121248 59200 121376
rect 880 120968 59120 121248
rect 880 120840 59200 120968
rect 880 120560 59120 120840
rect 880 120432 59200 120560
rect 880 120152 59120 120432
rect 880 120024 59200 120152
rect 880 119744 59120 120024
rect 880 119616 59200 119744
rect 880 119336 59120 119616
rect 880 119208 59200 119336
rect 880 118928 59120 119208
rect 880 118800 59200 118928
rect 880 118520 59120 118800
rect 880 118392 59200 118520
rect 880 118112 59120 118392
rect 880 117984 59200 118112
rect 880 117704 59120 117984
rect 880 117576 59200 117704
rect 880 117296 59120 117576
rect 880 117168 59200 117296
rect 880 116888 59120 117168
rect 880 116760 59200 116888
rect 880 116480 59120 116760
rect 880 116352 59200 116480
rect 880 116072 59120 116352
rect 880 115944 59200 116072
rect 880 115664 59120 115944
rect 880 115536 59200 115664
rect 880 115256 59120 115536
rect 880 115128 59200 115256
rect 880 114848 59120 115128
rect 880 114720 59200 114848
rect 880 114440 59120 114720
rect 880 114312 59200 114440
rect 880 114032 59120 114312
rect 880 113904 59200 114032
rect 880 113624 59120 113904
rect 880 113496 59200 113624
rect 880 113216 59120 113496
rect 880 113088 59200 113216
rect 880 112808 59120 113088
rect 880 112680 59200 112808
rect 880 112400 59120 112680
rect 880 112272 59200 112400
rect 880 111992 59120 112272
rect 880 111864 59200 111992
rect 880 111584 59120 111864
rect 880 111456 59200 111584
rect 880 111176 59120 111456
rect 880 111048 59200 111176
rect 880 110768 59120 111048
rect 880 110640 59200 110768
rect 880 110360 59120 110640
rect 880 110232 59200 110360
rect 880 109952 59120 110232
rect 880 109824 59200 109952
rect 880 109544 59120 109824
rect 880 109416 59200 109544
rect 880 109136 59120 109416
rect 880 109008 59200 109136
rect 880 108728 59120 109008
rect 880 108600 59200 108728
rect 880 108320 59120 108600
rect 880 108192 59200 108320
rect 880 107912 59120 108192
rect 880 107784 59200 107912
rect 880 107504 59120 107784
rect 880 107376 59200 107504
rect 880 107096 59120 107376
rect 880 106968 59200 107096
rect 880 106688 59120 106968
rect 880 106560 59200 106688
rect 880 106280 59120 106560
rect 880 106152 59200 106280
rect 880 105872 59120 106152
rect 880 105744 59200 105872
rect 880 105464 59120 105744
rect 880 105336 59200 105464
rect 880 105056 59120 105336
rect 880 104928 59200 105056
rect 880 104648 59120 104928
rect 880 104520 59200 104648
rect 880 104240 59120 104520
rect 880 104112 59200 104240
rect 880 103832 59120 104112
rect 880 103704 59200 103832
rect 880 103424 59120 103704
rect 880 103296 59200 103424
rect 880 103016 59120 103296
rect 880 102888 59200 103016
rect 880 102608 59120 102888
rect 880 102480 59200 102608
rect 880 102200 59120 102480
rect 880 102072 59200 102200
rect 880 101792 59120 102072
rect 880 101664 59200 101792
rect 880 101384 59120 101664
rect 880 101256 59200 101384
rect 880 100976 59120 101256
rect 880 100848 59200 100976
rect 880 100568 59120 100848
rect 880 100440 59200 100568
rect 880 100160 59120 100440
rect 880 100032 59200 100160
rect 880 99752 59120 100032
rect 880 99624 59200 99752
rect 880 99344 59120 99624
rect 880 99216 59200 99344
rect 880 98936 59120 99216
rect 880 98808 59200 98936
rect 880 98528 59120 98808
rect 880 98400 59200 98528
rect 880 98120 59120 98400
rect 880 97992 59200 98120
rect 880 97712 59120 97992
rect 880 97584 59200 97712
rect 880 97304 59120 97584
rect 880 97176 59200 97304
rect 880 96896 59120 97176
rect 880 96768 59200 96896
rect 880 96488 59120 96768
rect 880 96360 59200 96488
rect 880 96080 59120 96360
rect 880 95952 59200 96080
rect 880 95672 59120 95952
rect 880 95544 59200 95672
rect 880 95264 59120 95544
rect 880 95136 59200 95264
rect 880 94856 59120 95136
rect 880 94728 59200 94856
rect 880 94448 59120 94728
rect 880 94320 59200 94448
rect 880 94040 59120 94320
rect 880 93912 59200 94040
rect 880 93632 59120 93912
rect 880 93504 59200 93632
rect 880 93224 59120 93504
rect 880 93096 59200 93224
rect 880 92816 59120 93096
rect 880 92688 59200 92816
rect 880 92408 59120 92688
rect 880 92280 59200 92408
rect 880 92000 59120 92280
rect 880 91872 59200 92000
rect 880 91592 59120 91872
rect 880 91464 59200 91592
rect 880 91184 59120 91464
rect 880 91056 59200 91184
rect 880 90776 59120 91056
rect 880 90648 59200 90776
rect 880 90368 59120 90648
rect 880 90240 59200 90368
rect 880 89960 59120 90240
rect 880 89832 59200 89960
rect 880 89552 59120 89832
rect 880 89424 59200 89552
rect 880 89144 59120 89424
rect 880 89016 59200 89144
rect 880 88736 59120 89016
rect 880 88608 59200 88736
rect 880 88328 59120 88608
rect 880 88200 59200 88328
rect 880 87920 59120 88200
rect 880 87792 59200 87920
rect 880 87512 59120 87792
rect 880 87384 59200 87512
rect 880 87104 59120 87384
rect 880 86976 59200 87104
rect 880 86696 59120 86976
rect 880 86568 59200 86696
rect 880 86288 59120 86568
rect 880 86160 59200 86288
rect 880 85880 59120 86160
rect 880 85752 59200 85880
rect 880 85472 59120 85752
rect 880 85344 59200 85472
rect 880 85064 59120 85344
rect 880 84936 59200 85064
rect 880 84656 59120 84936
rect 880 84528 59200 84656
rect 880 84248 59120 84528
rect 880 84120 59200 84248
rect 880 83840 59120 84120
rect 880 83712 59200 83840
rect 880 83432 59120 83712
rect 880 83304 59200 83432
rect 880 83024 59120 83304
rect 880 82896 59200 83024
rect 880 82616 59120 82896
rect 880 82488 59200 82616
rect 880 82208 59120 82488
rect 880 82080 59200 82208
rect 880 81800 59120 82080
rect 880 81672 59200 81800
rect 880 81392 59120 81672
rect 880 81264 59200 81392
rect 880 80984 59120 81264
rect 880 80856 59200 80984
rect 880 80576 59120 80856
rect 880 80448 59200 80576
rect 880 80168 59120 80448
rect 880 80040 59200 80168
rect 880 79760 59120 80040
rect 880 79632 59200 79760
rect 880 79352 59120 79632
rect 880 79224 59200 79352
rect 880 78944 59120 79224
rect 880 78816 59200 78944
rect 880 78536 59120 78816
rect 880 78408 59200 78536
rect 880 78128 59120 78408
rect 880 78000 59200 78128
rect 880 77720 59120 78000
rect 880 77592 59200 77720
rect 880 77312 59120 77592
rect 880 77184 59200 77312
rect 880 76904 59120 77184
rect 880 76776 59200 76904
rect 880 76496 59120 76776
rect 880 76368 59200 76496
rect 880 76088 59120 76368
rect 880 75960 59200 76088
rect 880 75680 59120 75960
rect 880 75552 59200 75680
rect 880 75272 59120 75552
rect 880 75144 59200 75272
rect 880 74864 59120 75144
rect 880 74736 59200 74864
rect 880 74456 59120 74736
rect 880 74328 59200 74456
rect 880 74048 59120 74328
rect 880 73920 59200 74048
rect 880 73640 59120 73920
rect 880 73512 59200 73640
rect 880 73232 59120 73512
rect 880 73104 59200 73232
rect 880 72824 59120 73104
rect 880 72696 59200 72824
rect 880 72416 59120 72696
rect 880 72288 59200 72416
rect 880 72008 59120 72288
rect 880 71880 59200 72008
rect 880 71600 59120 71880
rect 880 71472 59200 71600
rect 880 71192 59120 71472
rect 880 71064 59200 71192
rect 880 70784 59120 71064
rect 880 70656 59200 70784
rect 880 70376 59120 70656
rect 880 70248 59200 70376
rect 880 69968 59120 70248
rect 880 69840 59200 69968
rect 880 69560 59120 69840
rect 880 69432 59200 69560
rect 880 69152 59120 69432
rect 880 69024 59200 69152
rect 880 68744 59120 69024
rect 880 68616 59200 68744
rect 880 68336 59120 68616
rect 880 68208 59200 68336
rect 880 67928 59120 68208
rect 880 67800 59200 67928
rect 880 67520 59120 67800
rect 880 67392 59200 67520
rect 880 67112 59120 67392
rect 880 66984 59200 67112
rect 880 66704 59120 66984
rect 880 66576 59200 66704
rect 880 66296 59120 66576
rect 880 66168 59200 66296
rect 880 65888 59120 66168
rect 880 65760 59200 65888
rect 880 65480 59120 65760
rect 880 65352 59200 65480
rect 880 65072 59120 65352
rect 880 64944 59200 65072
rect 880 64664 59120 64944
rect 880 64536 59200 64664
rect 880 64256 59120 64536
rect 880 64128 59200 64256
rect 880 63848 59120 64128
rect 880 63720 59200 63848
rect 880 63440 59120 63720
rect 880 63312 59200 63440
rect 880 63032 59120 63312
rect 880 62904 59200 63032
rect 880 62624 59120 62904
rect 880 62496 59200 62624
rect 880 62216 59120 62496
rect 880 62088 59200 62216
rect 880 61808 59120 62088
rect 880 61680 59200 61808
rect 880 61400 59120 61680
rect 880 61272 59200 61400
rect 880 60992 59120 61272
rect 880 60864 59200 60992
rect 880 60584 59120 60864
rect 880 60456 59200 60584
rect 880 60176 59120 60456
rect 880 60048 59200 60176
rect 880 59768 59120 60048
rect 880 59640 59200 59768
rect 880 59360 59120 59640
rect 880 59232 59200 59360
rect 880 58952 59120 59232
rect 880 58824 59200 58952
rect 880 58544 59120 58824
rect 880 58416 59200 58544
rect 880 58136 59120 58416
rect 880 58008 59200 58136
rect 880 57728 59120 58008
rect 880 57600 59200 57728
rect 880 57320 59120 57600
rect 880 57192 59200 57320
rect 880 56912 59120 57192
rect 880 56784 59200 56912
rect 880 56504 59120 56784
rect 880 56376 59200 56504
rect 880 56096 59120 56376
rect 880 55968 59200 56096
rect 880 55688 59120 55968
rect 880 55560 59200 55688
rect 880 55280 59120 55560
rect 880 55152 59200 55280
rect 880 54872 59120 55152
rect 880 54744 59200 54872
rect 880 54464 59120 54744
rect 880 54336 59200 54464
rect 880 54056 59120 54336
rect 880 53928 59200 54056
rect 880 53648 59120 53928
rect 880 53520 59200 53648
rect 880 53240 59120 53520
rect 880 53112 59200 53240
rect 880 52832 59120 53112
rect 880 52704 59200 52832
rect 880 52424 59120 52704
rect 880 52296 59200 52424
rect 880 52016 59120 52296
rect 880 51888 59200 52016
rect 880 51608 59120 51888
rect 880 51480 59200 51608
rect 880 51200 59120 51480
rect 880 51072 59200 51200
rect 880 50792 59120 51072
rect 880 50664 59200 50792
rect 880 50384 59120 50664
rect 880 50256 59200 50384
rect 880 49976 59120 50256
rect 880 49848 59200 49976
rect 880 49568 59120 49848
rect 880 49440 59200 49568
rect 880 49160 59120 49440
rect 880 49032 59200 49160
rect 880 48752 59120 49032
rect 880 48624 59200 48752
rect 880 48344 59120 48624
rect 880 48216 59200 48344
rect 880 47936 59120 48216
rect 880 47808 59200 47936
rect 880 47528 59120 47808
rect 880 47400 59200 47528
rect 880 47120 59120 47400
rect 880 46992 59200 47120
rect 880 46712 59120 46992
rect 880 46584 59200 46712
rect 880 46304 59120 46584
rect 880 46176 59200 46304
rect 880 45896 59120 46176
rect 880 45768 59200 45896
rect 880 45488 59120 45768
rect 880 45360 59200 45488
rect 880 45080 59120 45360
rect 880 44952 59200 45080
rect 880 44672 59120 44952
rect 880 44544 59200 44672
rect 880 44264 59120 44544
rect 880 44136 59200 44264
rect 880 43856 59120 44136
rect 880 43728 59200 43856
rect 880 43448 59120 43728
rect 880 43320 59200 43448
rect 880 43040 59120 43320
rect 880 42912 59200 43040
rect 880 42632 59120 42912
rect 880 42504 59200 42632
rect 880 42224 59120 42504
rect 880 42096 59200 42224
rect 880 41816 59120 42096
rect 880 41688 59200 41816
rect 880 41408 59120 41688
rect 880 41280 59200 41408
rect 880 41000 59120 41280
rect 880 40872 59200 41000
rect 880 40592 59120 40872
rect 880 40464 59200 40592
rect 880 40184 59120 40464
rect 880 40056 59200 40184
rect 880 39776 59120 40056
rect 880 39648 59200 39776
rect 880 39368 59120 39648
rect 880 39240 59200 39368
rect 880 38960 59120 39240
rect 880 38832 59200 38960
rect 880 38552 59120 38832
rect 880 38424 59200 38552
rect 880 38144 59120 38424
rect 880 38016 59200 38144
rect 880 37736 59120 38016
rect 880 37608 59200 37736
rect 880 37328 59120 37608
rect 880 37200 59200 37328
rect 880 36920 59120 37200
rect 880 36792 59200 36920
rect 880 36512 59120 36792
rect 880 36384 59200 36512
rect 880 36104 59120 36384
rect 880 35976 59200 36104
rect 880 35696 59120 35976
rect 880 35568 59200 35696
rect 880 35288 59120 35568
rect 880 35160 59200 35288
rect 880 34880 59120 35160
rect 880 34752 59200 34880
rect 880 34472 59120 34752
rect 880 34344 59200 34472
rect 880 34064 59120 34344
rect 880 33936 59200 34064
rect 880 33656 59120 33936
rect 880 33528 59200 33656
rect 880 33248 59120 33528
rect 880 33120 59200 33248
rect 880 32840 59120 33120
rect 880 32712 59200 32840
rect 880 32432 59120 32712
rect 880 32304 59200 32432
rect 880 32024 59120 32304
rect 880 31896 59200 32024
rect 880 31616 59120 31896
rect 880 31488 59200 31616
rect 880 31208 59120 31488
rect 880 31080 59200 31208
rect 880 30800 59120 31080
rect 880 30672 59200 30800
rect 880 30392 59120 30672
rect 880 30264 59200 30392
rect 880 29984 59120 30264
rect 880 29856 59200 29984
rect 880 29576 59120 29856
rect 880 29448 59200 29576
rect 880 29168 59120 29448
rect 880 29040 59200 29168
rect 880 28760 59120 29040
rect 880 28632 59200 28760
rect 880 28352 59120 28632
rect 880 28224 59200 28352
rect 880 27944 59120 28224
rect 880 27816 59200 27944
rect 880 27536 59120 27816
rect 880 27408 59200 27536
rect 880 27128 59120 27408
rect 880 27000 59200 27128
rect 880 26720 59120 27000
rect 880 26592 59200 26720
rect 880 26312 59120 26592
rect 880 26184 59200 26312
rect 880 25904 59120 26184
rect 880 25776 59200 25904
rect 880 25496 59120 25776
rect 880 25368 59200 25496
rect 880 25088 59120 25368
rect 880 24960 59200 25088
rect 880 24680 59120 24960
rect 880 24552 59200 24680
rect 880 24272 59120 24552
rect 880 24144 59200 24272
rect 880 23864 59120 24144
rect 880 23736 59200 23864
rect 880 23456 59120 23736
rect 880 23328 59200 23456
rect 880 23048 59120 23328
rect 880 22920 59200 23048
rect 880 22640 59120 22920
rect 880 22512 59200 22640
rect 880 22232 59120 22512
rect 800 22104 59200 22232
rect 800 21824 59120 22104
rect 800 21696 59200 21824
rect 800 21416 59120 21696
rect 800 21288 59200 21416
rect 800 21008 59120 21288
rect 800 20880 59200 21008
rect 800 20600 59120 20880
rect 800 20472 59200 20600
rect 800 20192 59120 20472
rect 800 20064 59200 20192
rect 800 19784 59120 20064
rect 800 19656 59200 19784
rect 800 19376 59120 19656
rect 800 19248 59200 19376
rect 800 18968 59120 19248
rect 800 18840 59200 18968
rect 800 18560 59120 18840
rect 800 18432 59200 18560
rect 800 18152 59120 18432
rect 800 18024 59200 18152
rect 800 17744 59120 18024
rect 800 17616 59200 17744
rect 800 17336 59120 17616
rect 800 17208 59200 17336
rect 800 16928 59120 17208
rect 800 16800 59200 16928
rect 800 16520 59120 16800
rect 800 16392 59200 16520
rect 800 16112 59120 16392
rect 800 15984 59200 16112
rect 800 15704 59120 15984
rect 800 2143 59200 15704
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
<< obsm4 >>
rect 430 2347 4128 151469
rect 4608 2347 19488 151469
rect 19968 2347 34848 151469
rect 35328 2347 50208 151469
rect 50688 2347 57717 151469
<< labels >>
rlabel metal3 s 0 22312 800 22432 6 c0_clk
port 1 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 c0_dbg_pc[0]
port 2 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 c0_dbg_pc[10]
port 3 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 c0_dbg_pc[11]
port 4 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 c0_dbg_pc[12]
port 5 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 c0_dbg_pc[13]
port 6 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 c0_dbg_pc[14]
port 7 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 c0_dbg_pc[15]
port 8 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 c0_dbg_pc[1]
port 9 nsew signal input
rlabel metal3 s 0 34280 800 34400 6 c0_dbg_pc[2]
port 10 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 c0_dbg_pc[3]
port 11 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 c0_dbg_pc[4]
port 12 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 c0_dbg_pc[5]
port 13 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 c0_dbg_pc[6]
port 14 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 c0_dbg_pc[7]
port 15 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 c0_dbg_pc[8]
port 16 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 c0_dbg_pc[9]
port 17 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 c0_dbg_r0[0]
port 18 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 c0_dbg_r0[10]
port 19 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 c0_dbg_r0[11]
port 20 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 c0_dbg_r0[12]
port 21 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 c0_dbg_r0[13]
port 22 nsew signal input
rlabel metal3 s 0 70456 800 70576 6 c0_dbg_r0[14]
port 23 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 c0_dbg_r0[15]
port 24 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 c0_dbg_r0[1]
port 25 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 c0_dbg_r0[2]
port 26 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 c0_dbg_r0[3]
port 27 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 c0_dbg_r0[4]
port 28 nsew signal input
rlabel metal3 s 0 44344 800 44464 6 c0_dbg_r0[5]
port 29 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 c0_dbg_r0[6]
port 30 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 c0_dbg_r0[7]
port 31 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 c0_dbg_r0[8]
port 32 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 c0_dbg_r0[9]
port 33 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 c0_disable
port 34 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 c0_i_core_int_sreg[0]
port 35 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 c0_i_core_int_sreg[10]
port 36 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 c0_i_core_int_sreg[11]
port 37 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 c0_i_core_int_sreg[12]
port 38 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 c0_i_core_int_sreg[13]
port 39 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 c0_i_core_int_sreg[14]
port 40 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 c0_i_core_int_sreg[15]
port 41 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 c0_i_core_int_sreg[1]
port 42 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 c0_i_core_int_sreg[2]
port 43 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 c0_i_core_int_sreg[3]
port 44 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 c0_i_core_int_sreg[4]
port 45 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 c0_i_core_int_sreg[5]
port 46 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 c0_i_core_int_sreg[6]
port 47 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 c0_i_core_int_sreg[7]
port 48 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 c0_i_core_int_sreg[8]
port 49 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 c0_i_core_int_sreg[9]
port 50 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 c0_i_irq
port 51 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 c0_i_mc_core_int
port 52 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 c0_i_mem_ack
port 53 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 c0_i_mem_data[0]
port 54 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 c0_i_mem_data[10]
port 55 nsew signal output
rlabel metal3 s 0 62840 800 62960 6 c0_i_mem_data[11]
port 56 nsew signal output
rlabel metal3 s 0 65560 800 65680 6 c0_i_mem_data[12]
port 57 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 c0_i_mem_data[13]
port 58 nsew signal output
rlabel metal3 s 0 71000 800 71120 6 c0_i_mem_data[14]
port 59 nsew signal output
rlabel metal3 s 0 73720 800 73840 6 c0_i_mem_data[15]
port 60 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 c0_i_mem_data[1]
port 61 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 c0_i_mem_data[2]
port 62 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 c0_i_mem_data[3]
port 63 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 c0_i_mem_data[4]
port 64 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 c0_i_mem_data[5]
port 65 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 c0_i_mem_data[6]
port 66 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 c0_i_mem_data[7]
port 67 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 c0_i_mem_data[8]
port 68 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 c0_i_mem_data[9]
port 69 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 c0_i_mem_exception
port 70 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 c0_i_req_data[0]
port 71 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 c0_i_req_data[10]
port 72 nsew signal output
rlabel metal3 s 0 63112 800 63232 6 c0_i_req_data[11]
port 73 nsew signal output
rlabel metal3 s 0 65832 800 65952 6 c0_i_req_data[12]
port 74 nsew signal output
rlabel metal3 s 0 68552 800 68672 6 c0_i_req_data[13]
port 75 nsew signal output
rlabel metal3 s 0 71272 800 71392 6 c0_i_req_data[14]
port 76 nsew signal output
rlabel metal3 s 0 73992 800 74112 6 c0_i_req_data[15]
port 77 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 c0_i_req_data[16]
port 78 nsew signal output
rlabel metal3 s 0 75896 800 76016 6 c0_i_req_data[17]
port 79 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 c0_i_req_data[18]
port 80 nsew signal output
rlabel metal3 s 0 76440 800 76560 6 c0_i_req_data[19]
port 81 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 c0_i_req_data[1]
port 82 nsew signal output
rlabel metal3 s 0 76712 800 76832 6 c0_i_req_data[20]
port 83 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 c0_i_req_data[21]
port 84 nsew signal output
rlabel metal3 s 0 77256 800 77376 6 c0_i_req_data[22]
port 85 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 c0_i_req_data[23]
port 86 nsew signal output
rlabel metal3 s 0 77800 800 77920 6 c0_i_req_data[24]
port 87 nsew signal output
rlabel metal3 s 0 78072 800 78192 6 c0_i_req_data[25]
port 88 nsew signal output
rlabel metal3 s 0 78344 800 78464 6 c0_i_req_data[26]
port 89 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 c0_i_req_data[27]
port 90 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 c0_i_req_data[28]
port 91 nsew signal output
rlabel metal3 s 0 79160 800 79280 6 c0_i_req_data[29]
port 92 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 c0_i_req_data[2]
port 93 nsew signal output
rlabel metal3 s 0 79432 800 79552 6 c0_i_req_data[30]
port 94 nsew signal output
rlabel metal3 s 0 79704 800 79824 6 c0_i_req_data[31]
port 95 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 c0_i_req_data[3]
port 96 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 c0_i_req_data[4]
port 97 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 c0_i_req_data[5]
port 98 nsew signal output
rlabel metal3 s 0 48424 800 48544 6 c0_i_req_data[6]
port 99 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 c0_i_req_data[7]
port 100 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 c0_i_req_data[8]
port 101 nsew signal output
rlabel metal3 s 0 57672 800 57792 6 c0_i_req_data[9]
port 102 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 c0_i_req_data_valid
port 103 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 c0_o_c_data_page
port 104 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 c0_o_c_instr_long
port 105 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 c0_o_c_instr_page
port 106 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 c0_o_icache_flush
port 107 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 c0_o_instr_long_addr[0]
port 108 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 c0_o_instr_long_addr[1]
port 109 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 c0_o_instr_long_addr[2]
port 110 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 c0_o_instr_long_addr[3]
port 111 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 c0_o_instr_long_addr[4]
port 112 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 c0_o_instr_long_addr[5]
port 113 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 c0_o_instr_long_addr[6]
port 114 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 c0_o_instr_long_addr[7]
port 115 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 c0_o_mem_addr[0]
port 116 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 c0_o_mem_addr[10]
port 117 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 c0_o_mem_addr[11]
port 118 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 c0_o_mem_addr[12]
port 119 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 c0_o_mem_addr[13]
port 120 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 c0_o_mem_addr[14]
port 121 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 c0_o_mem_addr[15]
port 122 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 c0_o_mem_addr[1]
port 123 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 c0_o_mem_addr[2]
port 124 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 c0_o_mem_addr[3]
port 125 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 c0_o_mem_addr[4]
port 126 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 c0_o_mem_addr[5]
port 127 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 c0_o_mem_addr[6]
port 128 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 c0_o_mem_addr[7]
port 129 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 c0_o_mem_addr[8]
port 130 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 c0_o_mem_addr[9]
port 131 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 c0_o_mem_data[0]
port 132 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 c0_o_mem_data[10]
port 133 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 c0_o_mem_data[11]
port 134 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 c0_o_mem_data[12]
port 135 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 c0_o_mem_data[13]
port 136 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 c0_o_mem_data[14]
port 137 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 c0_o_mem_data[15]
port 138 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 c0_o_mem_data[1]
port 139 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 c0_o_mem_data[2]
port 140 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 c0_o_mem_data[3]
port 141 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 c0_o_mem_data[4]
port 142 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 c0_o_mem_data[5]
port 143 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 c0_o_mem_data[6]
port 144 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 c0_o_mem_data[7]
port 145 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 c0_o_mem_data[8]
port 146 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 c0_o_mem_data[9]
port 147 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 c0_o_mem_high_addr[0]
port 148 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 c0_o_mem_high_addr[1]
port 149 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 c0_o_mem_high_addr[2]
port 150 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 c0_o_mem_high_addr[3]
port 151 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 c0_o_mem_high_addr[4]
port 152 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 c0_o_mem_high_addr[5]
port 153 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 c0_o_mem_high_addr[6]
port 154 nsew signal input
rlabel metal3 s 0 52776 800 52896 6 c0_o_mem_high_addr[7]
port 155 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 c0_o_mem_long_mode
port 156 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 c0_o_mem_req
port 157 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 c0_o_mem_sel[0]
port 158 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 c0_o_mem_sel[1]
port 159 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 c0_o_mem_we
port 160 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 c0_o_req_active
port 161 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 c0_o_req_addr[0]
port 162 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 c0_o_req_addr[10]
port 163 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 c0_o_req_addr[11]
port 164 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 c0_o_req_addr[12]
port 165 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 c0_o_req_addr[13]
port 166 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 c0_o_req_addr[14]
port 167 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 c0_o_req_addr[15]
port 168 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 c0_o_req_addr[1]
port 169 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 c0_o_req_addr[2]
port 170 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 c0_o_req_addr[3]
port 171 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 c0_o_req_addr[4]
port 172 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 c0_o_req_addr[5]
port 173 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 c0_o_req_addr[6]
port 174 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 c0_o_req_addr[7]
port 175 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 c0_o_req_addr[8]
port 176 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 c0_o_req_addr[9]
port 177 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 c0_o_req_ppl_submit
port 178 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 c0_rst
port 179 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 c0_sr_bus_addr[0]
port 180 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 c0_sr_bus_addr[10]
port 181 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 c0_sr_bus_addr[11]
port 182 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 c0_sr_bus_addr[12]
port 183 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 c0_sr_bus_addr[13]
port 184 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 c0_sr_bus_addr[14]
port 185 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 c0_sr_bus_addr[15]
port 186 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 c0_sr_bus_addr[1]
port 187 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 c0_sr_bus_addr[2]
port 188 nsew signal input
rlabel metal3 s 0 40264 800 40384 6 c0_sr_bus_addr[3]
port 189 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 c0_sr_bus_addr[4]
port 190 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 c0_sr_bus_addr[5]
port 191 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 c0_sr_bus_addr[6]
port 192 nsew signal input
rlabel metal3 s 0 53320 800 53440 6 c0_sr_bus_addr[7]
port 193 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 c0_sr_bus_addr[8]
port 194 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 c0_sr_bus_addr[9]
port 195 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 c0_sr_bus_data_o[0]
port 196 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 c0_sr_bus_data_o[10]
port 197 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 c0_sr_bus_data_o[11]
port 198 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 c0_sr_bus_data_o[12]
port 199 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 c0_sr_bus_data_o[13]
port 200 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 c0_sr_bus_data_o[14]
port 201 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 c0_sr_bus_data_o[15]
port 202 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 c0_sr_bus_data_o[1]
port 203 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 c0_sr_bus_data_o[2]
port 204 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 c0_sr_bus_data_o[3]
port 205 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 c0_sr_bus_data_o[4]
port 206 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 c0_sr_bus_data_o[5]
port 207 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 c0_sr_bus_data_o[6]
port 208 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 c0_sr_bus_data_o[7]
port 209 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 c0_sr_bus_data_o[8]
port 210 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 c0_sr_bus_data_o[9]
port 211 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 c0_sr_bus_we
port 212 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 c1_clk
port 213 nsew signal output
rlabel metal3 s 0 84872 800 84992 6 c1_dbg_pc[0]
port 214 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 c1_dbg_pc[10]
port 215 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 c1_dbg_pc[11]
port 216 nsew signal input
rlabel metal3 s 0 122408 800 122528 6 c1_dbg_pc[12]
port 217 nsew signal input
rlabel metal3 s 0 125128 800 125248 6 c1_dbg_pc[13]
port 218 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 c1_dbg_pc[14]
port 219 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 c1_dbg_pc[15]
port 220 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 c1_dbg_pc[1]
port 221 nsew signal input
rlabel metal3 s 0 91944 800 92064 6 c1_dbg_pc[2]
port 222 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 c1_dbg_pc[3]
port 223 nsew signal input
rlabel metal3 s 0 98472 800 98592 6 c1_dbg_pc[4]
port 224 nsew signal input
rlabel metal3 s 0 101736 800 101856 6 c1_dbg_pc[5]
port 225 nsew signal input
rlabel metal3 s 0 105000 800 105120 6 c1_dbg_pc[6]
port 226 nsew signal input
rlabel metal3 s 0 108264 800 108384 6 c1_dbg_pc[7]
port 227 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 c1_dbg_pc[8]
port 228 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 c1_dbg_pc[9]
port 229 nsew signal input
rlabel metal3 s 0 85144 800 85264 6 c1_dbg_r0[0]
port 230 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 c1_dbg_r0[10]
port 231 nsew signal input
rlabel metal3 s 0 119960 800 120080 6 c1_dbg_r0[11]
port 232 nsew signal input
rlabel metal3 s 0 122680 800 122800 6 c1_dbg_r0[12]
port 233 nsew signal input
rlabel metal3 s 0 125400 800 125520 6 c1_dbg_r0[13]
port 234 nsew signal input
rlabel metal3 s 0 128120 800 128240 6 c1_dbg_r0[14]
port 235 nsew signal input
rlabel metal3 s 0 130840 800 130960 6 c1_dbg_r0[15]
port 236 nsew signal input
rlabel metal3 s 0 88680 800 88800 6 c1_dbg_r0[1]
port 237 nsew signal input
rlabel metal3 s 0 92216 800 92336 6 c1_dbg_r0[2]
port 238 nsew signal input
rlabel metal3 s 0 95480 800 95600 6 c1_dbg_r0[3]
port 239 nsew signal input
rlabel metal3 s 0 98744 800 98864 6 c1_dbg_r0[4]
port 240 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 c1_dbg_r0[5]
port 241 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 c1_dbg_r0[6]
port 242 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 c1_dbg_r0[7]
port 243 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 c1_dbg_r0[8]
port 244 nsew signal input
rlabel metal3 s 0 114520 800 114640 6 c1_dbg_r0[9]
port 245 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 c1_disable
port 246 nsew signal output
rlabel metal3 s 0 85416 800 85536 6 c1_i_core_int_sreg[0]
port 247 nsew signal output
rlabel metal3 s 0 117512 800 117632 6 c1_i_core_int_sreg[10]
port 248 nsew signal output
rlabel metal3 s 0 120232 800 120352 6 c1_i_core_int_sreg[11]
port 249 nsew signal output
rlabel metal3 s 0 122952 800 123072 6 c1_i_core_int_sreg[12]
port 250 nsew signal output
rlabel metal3 s 0 125672 800 125792 6 c1_i_core_int_sreg[13]
port 251 nsew signal output
rlabel metal3 s 0 128392 800 128512 6 c1_i_core_int_sreg[14]
port 252 nsew signal output
rlabel metal3 s 0 131112 800 131232 6 c1_i_core_int_sreg[15]
port 253 nsew signal output
rlabel metal3 s 0 88952 800 89072 6 c1_i_core_int_sreg[1]
port 254 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 c1_i_core_int_sreg[2]
port 255 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 c1_i_core_int_sreg[3]
port 256 nsew signal output
rlabel metal3 s 0 99016 800 99136 6 c1_i_core_int_sreg[4]
port 257 nsew signal output
rlabel metal3 s 0 102280 800 102400 6 c1_i_core_int_sreg[5]
port 258 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 c1_i_core_int_sreg[6]
port 259 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 c1_i_core_int_sreg[7]
port 260 nsew signal output
rlabel metal3 s 0 112072 800 112192 6 c1_i_core_int_sreg[8]
port 261 nsew signal output
rlabel metal3 s 0 114792 800 114912 6 c1_i_core_int_sreg[9]
port 262 nsew signal output
rlabel metal3 s 0 80520 800 80640 6 c1_i_irq
port 263 nsew signal output
rlabel metal3 s 0 80792 800 80912 6 c1_i_mc_core_int
port 264 nsew signal output
rlabel metal3 s 0 81064 800 81184 6 c1_i_mem_ack
port 265 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 c1_i_mem_data[0]
port 266 nsew signal output
rlabel metal3 s 0 117784 800 117904 6 c1_i_mem_data[10]
port 267 nsew signal output
rlabel metal3 s 0 120504 800 120624 6 c1_i_mem_data[11]
port 268 nsew signal output
rlabel metal3 s 0 123224 800 123344 6 c1_i_mem_data[12]
port 269 nsew signal output
rlabel metal3 s 0 125944 800 126064 6 c1_i_mem_data[13]
port 270 nsew signal output
rlabel metal3 s 0 128664 800 128784 6 c1_i_mem_data[14]
port 271 nsew signal output
rlabel metal3 s 0 131384 800 131504 6 c1_i_mem_data[15]
port 272 nsew signal output
rlabel metal3 s 0 89224 800 89344 6 c1_i_mem_data[1]
port 273 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 c1_i_mem_data[2]
port 274 nsew signal output
rlabel metal3 s 0 96024 800 96144 6 c1_i_mem_data[3]
port 275 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 c1_i_mem_data[4]
port 276 nsew signal output
rlabel metal3 s 0 102552 800 102672 6 c1_i_mem_data[5]
port 277 nsew signal output
rlabel metal3 s 0 105816 800 105936 6 c1_i_mem_data[6]
port 278 nsew signal output
rlabel metal3 s 0 109080 800 109200 6 c1_i_mem_data[7]
port 279 nsew signal output
rlabel metal3 s 0 112344 800 112464 6 c1_i_mem_data[8]
port 280 nsew signal output
rlabel metal3 s 0 115064 800 115184 6 c1_i_mem_data[9]
port 281 nsew signal output
rlabel metal3 s 0 81336 800 81456 6 c1_i_mem_exception
port 282 nsew signal output
rlabel metal3 s 0 85960 800 86080 6 c1_i_req_data[0]
port 283 nsew signal output
rlabel metal3 s 0 118056 800 118176 6 c1_i_req_data[10]
port 284 nsew signal output
rlabel metal3 s 0 120776 800 120896 6 c1_i_req_data[11]
port 285 nsew signal output
rlabel metal3 s 0 123496 800 123616 6 c1_i_req_data[12]
port 286 nsew signal output
rlabel metal3 s 0 126216 800 126336 6 c1_i_req_data[13]
port 287 nsew signal output
rlabel metal3 s 0 128936 800 129056 6 c1_i_req_data[14]
port 288 nsew signal output
rlabel metal3 s 0 131656 800 131776 6 c1_i_req_data[15]
port 289 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 c1_i_req_data[16]
port 290 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 c1_i_req_data[17]
port 291 nsew signal output
rlabel metal3 s 0 133832 800 133952 6 c1_i_req_data[18]
port 292 nsew signal output
rlabel metal3 s 0 134104 800 134224 6 c1_i_req_data[19]
port 293 nsew signal output
rlabel metal3 s 0 89496 800 89616 6 c1_i_req_data[1]
port 294 nsew signal output
rlabel metal3 s 0 134376 800 134496 6 c1_i_req_data[20]
port 295 nsew signal output
rlabel metal3 s 0 134648 800 134768 6 c1_i_req_data[21]
port 296 nsew signal output
rlabel metal3 s 0 134920 800 135040 6 c1_i_req_data[22]
port 297 nsew signal output
rlabel metal3 s 0 135192 800 135312 6 c1_i_req_data[23]
port 298 nsew signal output
rlabel metal3 s 0 135464 800 135584 6 c1_i_req_data[24]
port 299 nsew signal output
rlabel metal3 s 0 135736 800 135856 6 c1_i_req_data[25]
port 300 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 c1_i_req_data[26]
port 301 nsew signal output
rlabel metal3 s 0 136280 800 136400 6 c1_i_req_data[27]
port 302 nsew signal output
rlabel metal3 s 0 136552 800 136672 6 c1_i_req_data[28]
port 303 nsew signal output
rlabel metal3 s 0 136824 800 136944 6 c1_i_req_data[29]
port 304 nsew signal output
rlabel metal3 s 0 93032 800 93152 6 c1_i_req_data[2]
port 305 nsew signal output
rlabel metal3 s 0 137096 800 137216 6 c1_i_req_data[30]
port 306 nsew signal output
rlabel metal3 s 0 137368 800 137488 6 c1_i_req_data[31]
port 307 nsew signal output
rlabel metal3 s 0 96296 800 96416 6 c1_i_req_data[3]
port 308 nsew signal output
rlabel metal3 s 0 99560 800 99680 6 c1_i_req_data[4]
port 309 nsew signal output
rlabel metal3 s 0 102824 800 102944 6 c1_i_req_data[5]
port 310 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 c1_i_req_data[6]
port 311 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 c1_i_req_data[7]
port 312 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 c1_i_req_data[8]
port 313 nsew signal output
rlabel metal3 s 0 115336 800 115456 6 c1_i_req_data[9]
port 314 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 c1_i_req_data_valid
port 315 nsew signal output
rlabel metal3 s 0 81880 800 82000 6 c1_o_c_data_page
port 316 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 c1_o_c_instr_long
port 317 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 c1_o_c_instr_page
port 318 nsew signal input
rlabel metal3 s 0 82696 800 82816 6 c1_o_icache_flush
port 319 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 c1_o_instr_long_addr[0]
port 320 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 c1_o_instr_long_addr[1]
port 321 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 c1_o_instr_long_addr[2]
port 322 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 c1_o_instr_long_addr[3]
port 323 nsew signal input
rlabel metal3 s 0 99832 800 99952 6 c1_o_instr_long_addr[4]
port 324 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 c1_o_instr_long_addr[5]
port 325 nsew signal input
rlabel metal3 s 0 106360 800 106480 6 c1_o_instr_long_addr[6]
port 326 nsew signal input
rlabel metal3 s 0 109624 800 109744 6 c1_o_instr_long_addr[7]
port 327 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 c1_o_mem_addr[0]
port 328 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 c1_o_mem_addr[10]
port 329 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 c1_o_mem_addr[11]
port 330 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 c1_o_mem_addr[12]
port 331 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 c1_o_mem_addr[13]
port 332 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 c1_o_mem_addr[14]
port 333 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 c1_o_mem_addr[15]
port 334 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 c1_o_mem_addr[1]
port 335 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 c1_o_mem_addr[2]
port 336 nsew signal input
rlabel metal3 s 0 96840 800 96960 6 c1_o_mem_addr[3]
port 337 nsew signal input
rlabel metal3 s 0 100104 800 100224 6 c1_o_mem_addr[4]
port 338 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 c1_o_mem_addr[5]
port 339 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 c1_o_mem_addr[6]
port 340 nsew signal input
rlabel metal3 s 0 109896 800 110016 6 c1_o_mem_addr[7]
port 341 nsew signal input
rlabel metal3 s 0 112888 800 113008 6 c1_o_mem_addr[8]
port 342 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 c1_o_mem_addr[9]
port 343 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 c1_o_mem_data[0]
port 344 nsew signal input
rlabel metal3 s 0 118600 800 118720 6 c1_o_mem_data[10]
port 345 nsew signal input
rlabel metal3 s 0 121320 800 121440 6 c1_o_mem_data[11]
port 346 nsew signal input
rlabel metal3 s 0 124040 800 124160 6 c1_o_mem_data[12]
port 347 nsew signal input
rlabel metal3 s 0 126760 800 126880 6 c1_o_mem_data[13]
port 348 nsew signal input
rlabel metal3 s 0 129480 800 129600 6 c1_o_mem_data[14]
port 349 nsew signal input
rlabel metal3 s 0 132200 800 132320 6 c1_o_mem_data[15]
port 350 nsew signal input
rlabel metal3 s 0 90312 800 90432 6 c1_o_mem_data[1]
port 351 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 c1_o_mem_data[2]
port 352 nsew signal input
rlabel metal3 s 0 97112 800 97232 6 c1_o_mem_data[3]
port 353 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 c1_o_mem_data[4]
port 354 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 c1_o_mem_data[5]
port 355 nsew signal input
rlabel metal3 s 0 106904 800 107024 6 c1_o_mem_data[6]
port 356 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 c1_o_mem_data[7]
port 357 nsew signal input
rlabel metal3 s 0 113160 800 113280 6 c1_o_mem_data[8]
port 358 nsew signal input
rlabel metal3 s 0 115880 800 116000 6 c1_o_mem_data[9]
port 359 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 c1_o_mem_high_addr[0]
port 360 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 c1_o_mem_high_addr[1]
port 361 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 c1_o_mem_high_addr[2]
port 362 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 c1_o_mem_high_addr[3]
port 363 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 c1_o_mem_high_addr[4]
port 364 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 c1_o_mem_high_addr[5]
port 365 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 c1_o_mem_high_addr[6]
port 366 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 c1_o_mem_high_addr[7]
port 367 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 c1_o_mem_long_mode
port 368 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 c1_o_mem_req
port 369 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 c1_o_mem_sel[0]
port 370 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 c1_o_mem_sel[1]
port 371 nsew signal input
rlabel metal3 s 0 83512 800 83632 6 c1_o_mem_we
port 372 nsew signal input
rlabel metal3 s 0 83784 800 83904 6 c1_o_req_active
port 373 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 c1_o_req_addr[0]
port 374 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 c1_o_req_addr[10]
port 375 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 c1_o_req_addr[11]
port 376 nsew signal input
rlabel metal3 s 0 124312 800 124432 6 c1_o_req_addr[12]
port 377 nsew signal input
rlabel metal3 s 0 127032 800 127152 6 c1_o_req_addr[13]
port 378 nsew signal input
rlabel metal3 s 0 129752 800 129872 6 c1_o_req_addr[14]
port 379 nsew signal input
rlabel metal3 s 0 132472 800 132592 6 c1_o_req_addr[15]
port 380 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 c1_o_req_addr[1]
port 381 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 c1_o_req_addr[2]
port 382 nsew signal input
rlabel metal3 s 0 97656 800 97776 6 c1_o_req_addr[3]
port 383 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 c1_o_req_addr[4]
port 384 nsew signal input
rlabel metal3 s 0 104184 800 104304 6 c1_o_req_addr[5]
port 385 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 c1_o_req_addr[6]
port 386 nsew signal input
rlabel metal3 s 0 110712 800 110832 6 c1_o_req_addr[7]
port 387 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 c1_o_req_addr[8]
port 388 nsew signal input
rlabel metal3 s 0 116152 800 116272 6 c1_o_req_addr[9]
port 389 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 c1_o_req_ppl_submit
port 390 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 c1_rst
port 391 nsew signal output
rlabel metal3 s 0 87864 800 87984 6 c1_sr_bus_addr[0]
port 392 nsew signal input
rlabel metal3 s 0 119144 800 119264 6 c1_sr_bus_addr[10]
port 393 nsew signal input
rlabel metal3 s 0 121864 800 121984 6 c1_sr_bus_addr[11]
port 394 nsew signal input
rlabel metal3 s 0 124584 800 124704 6 c1_sr_bus_addr[12]
port 395 nsew signal input
rlabel metal3 s 0 127304 800 127424 6 c1_sr_bus_addr[13]
port 396 nsew signal input
rlabel metal3 s 0 130024 800 130144 6 c1_sr_bus_addr[14]
port 397 nsew signal input
rlabel metal3 s 0 132744 800 132864 6 c1_sr_bus_addr[15]
port 398 nsew signal input
rlabel metal3 s 0 91400 800 91520 6 c1_sr_bus_addr[1]
port 399 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 c1_sr_bus_addr[2]
port 400 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 c1_sr_bus_addr[3]
port 401 nsew signal input
rlabel metal3 s 0 101192 800 101312 6 c1_sr_bus_addr[4]
port 402 nsew signal input
rlabel metal3 s 0 104456 800 104576 6 c1_sr_bus_addr[5]
port 403 nsew signal input
rlabel metal3 s 0 107720 800 107840 6 c1_sr_bus_addr[6]
port 404 nsew signal input
rlabel metal3 s 0 110984 800 111104 6 c1_sr_bus_addr[7]
port 405 nsew signal input
rlabel metal3 s 0 113704 800 113824 6 c1_sr_bus_addr[8]
port 406 nsew signal input
rlabel metal3 s 0 116424 800 116544 6 c1_sr_bus_addr[9]
port 407 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 c1_sr_bus_data_o[0]
port 408 nsew signal input
rlabel metal3 s 0 119416 800 119536 6 c1_sr_bus_data_o[10]
port 409 nsew signal input
rlabel metal3 s 0 122136 800 122256 6 c1_sr_bus_data_o[11]
port 410 nsew signal input
rlabel metal3 s 0 124856 800 124976 6 c1_sr_bus_data_o[12]
port 411 nsew signal input
rlabel metal3 s 0 127576 800 127696 6 c1_sr_bus_data_o[13]
port 412 nsew signal input
rlabel metal3 s 0 130296 800 130416 6 c1_sr_bus_data_o[14]
port 413 nsew signal input
rlabel metal3 s 0 133016 800 133136 6 c1_sr_bus_data_o[15]
port 414 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 c1_sr_bus_data_o[1]
port 415 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 c1_sr_bus_data_o[2]
port 416 nsew signal input
rlabel metal3 s 0 98200 800 98320 6 c1_sr_bus_data_o[3]
port 417 nsew signal input
rlabel metal3 s 0 101464 800 101584 6 c1_sr_bus_data_o[4]
port 418 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 c1_sr_bus_data_o[5]
port 419 nsew signal input
rlabel metal3 s 0 107992 800 108112 6 c1_sr_bus_data_o[6]
port 420 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 c1_sr_bus_data_o[7]
port 421 nsew signal input
rlabel metal3 s 0 113976 800 114096 6 c1_sr_bus_data_o[8]
port 422 nsew signal input
rlabel metal3 s 0 116696 800 116816 6 c1_sr_bus_data_o[9]
port 423 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 c1_sr_bus_we
port 424 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 core_clock
port 425 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 core_reset
port 426 nsew signal input
rlabel metal3 s 59200 15784 60000 15904 6 dcache_clk
port 427 nsew signal output
rlabel metal3 s 59200 16192 60000 16312 6 dcache_mem_ack
port 428 nsew signal input
rlabel metal3 s 59200 21088 60000 21208 6 dcache_mem_addr[0]
port 429 nsew signal output
rlabel metal3 s 59200 47200 60000 47320 6 dcache_mem_addr[10]
port 430 nsew signal output
rlabel metal3 s 59200 49648 60000 49768 6 dcache_mem_addr[11]
port 431 nsew signal output
rlabel metal3 s 59200 52096 60000 52216 6 dcache_mem_addr[12]
port 432 nsew signal output
rlabel metal3 s 59200 54544 60000 54664 6 dcache_mem_addr[13]
port 433 nsew signal output
rlabel metal3 s 59200 56992 60000 57112 6 dcache_mem_addr[14]
port 434 nsew signal output
rlabel metal3 s 59200 59440 60000 59560 6 dcache_mem_addr[15]
port 435 nsew signal output
rlabel metal3 s 59200 61888 60000 62008 6 dcache_mem_addr[16]
port 436 nsew signal output
rlabel metal3 s 59200 62704 60000 62824 6 dcache_mem_addr[17]
port 437 nsew signal output
rlabel metal3 s 59200 63520 60000 63640 6 dcache_mem_addr[18]
port 438 nsew signal output
rlabel metal3 s 59200 64336 60000 64456 6 dcache_mem_addr[19]
port 439 nsew signal output
rlabel metal3 s 59200 24352 60000 24472 6 dcache_mem_addr[1]
port 440 nsew signal output
rlabel metal3 s 59200 65152 60000 65272 6 dcache_mem_addr[20]
port 441 nsew signal output
rlabel metal3 s 59200 65968 60000 66088 6 dcache_mem_addr[21]
port 442 nsew signal output
rlabel metal3 s 59200 66784 60000 66904 6 dcache_mem_addr[22]
port 443 nsew signal output
rlabel metal3 s 59200 67600 60000 67720 6 dcache_mem_addr[23]
port 444 nsew signal output
rlabel metal3 s 59200 27616 60000 27736 6 dcache_mem_addr[2]
port 445 nsew signal output
rlabel metal3 s 59200 30064 60000 30184 6 dcache_mem_addr[3]
port 446 nsew signal output
rlabel metal3 s 59200 32512 60000 32632 6 dcache_mem_addr[4]
port 447 nsew signal output
rlabel metal3 s 59200 34960 60000 35080 6 dcache_mem_addr[5]
port 448 nsew signal output
rlabel metal3 s 59200 37408 60000 37528 6 dcache_mem_addr[6]
port 449 nsew signal output
rlabel metal3 s 59200 39856 60000 39976 6 dcache_mem_addr[7]
port 450 nsew signal output
rlabel metal3 s 59200 42304 60000 42424 6 dcache_mem_addr[8]
port 451 nsew signal output
rlabel metal3 s 59200 44752 60000 44872 6 dcache_mem_addr[9]
port 452 nsew signal output
rlabel metal3 s 59200 16600 60000 16720 6 dcache_mem_cache_enable
port 453 nsew signal output
rlabel metal3 s 59200 17008 60000 17128 6 dcache_mem_exception
port 454 nsew signal input
rlabel metal3 s 59200 21496 60000 21616 6 dcache_mem_i_data[0]
port 455 nsew signal output
rlabel metal3 s 59200 47608 60000 47728 6 dcache_mem_i_data[10]
port 456 nsew signal output
rlabel metal3 s 59200 50056 60000 50176 6 dcache_mem_i_data[11]
port 457 nsew signal output
rlabel metal3 s 59200 52504 60000 52624 6 dcache_mem_i_data[12]
port 458 nsew signal output
rlabel metal3 s 59200 54952 60000 55072 6 dcache_mem_i_data[13]
port 459 nsew signal output
rlabel metal3 s 59200 57400 60000 57520 6 dcache_mem_i_data[14]
port 460 nsew signal output
rlabel metal3 s 59200 59848 60000 59968 6 dcache_mem_i_data[15]
port 461 nsew signal output
rlabel metal3 s 59200 24760 60000 24880 6 dcache_mem_i_data[1]
port 462 nsew signal output
rlabel metal3 s 59200 28024 60000 28144 6 dcache_mem_i_data[2]
port 463 nsew signal output
rlabel metal3 s 59200 30472 60000 30592 6 dcache_mem_i_data[3]
port 464 nsew signal output
rlabel metal3 s 59200 32920 60000 33040 6 dcache_mem_i_data[4]
port 465 nsew signal output
rlabel metal3 s 59200 35368 60000 35488 6 dcache_mem_i_data[5]
port 466 nsew signal output
rlabel metal3 s 59200 37816 60000 37936 6 dcache_mem_i_data[6]
port 467 nsew signal output
rlabel metal3 s 59200 40264 60000 40384 6 dcache_mem_i_data[7]
port 468 nsew signal output
rlabel metal3 s 59200 42712 60000 42832 6 dcache_mem_i_data[8]
port 469 nsew signal output
rlabel metal3 s 59200 45160 60000 45280 6 dcache_mem_i_data[9]
port 470 nsew signal output
rlabel metal3 s 59200 21904 60000 22024 6 dcache_mem_o_data[0]
port 471 nsew signal input
rlabel metal3 s 59200 48016 60000 48136 6 dcache_mem_o_data[10]
port 472 nsew signal input
rlabel metal3 s 59200 50464 60000 50584 6 dcache_mem_o_data[11]
port 473 nsew signal input
rlabel metal3 s 59200 52912 60000 53032 6 dcache_mem_o_data[12]
port 474 nsew signal input
rlabel metal3 s 59200 55360 60000 55480 6 dcache_mem_o_data[13]
port 475 nsew signal input
rlabel metal3 s 59200 57808 60000 57928 6 dcache_mem_o_data[14]
port 476 nsew signal input
rlabel metal3 s 59200 60256 60000 60376 6 dcache_mem_o_data[15]
port 477 nsew signal input
rlabel metal3 s 59200 25168 60000 25288 6 dcache_mem_o_data[1]
port 478 nsew signal input
rlabel metal3 s 59200 28432 60000 28552 6 dcache_mem_o_data[2]
port 479 nsew signal input
rlabel metal3 s 59200 30880 60000 31000 6 dcache_mem_o_data[3]
port 480 nsew signal input
rlabel metal3 s 59200 33328 60000 33448 6 dcache_mem_o_data[4]
port 481 nsew signal input
rlabel metal3 s 59200 35776 60000 35896 6 dcache_mem_o_data[5]
port 482 nsew signal input
rlabel metal3 s 59200 38224 60000 38344 6 dcache_mem_o_data[6]
port 483 nsew signal input
rlabel metal3 s 59200 40672 60000 40792 6 dcache_mem_o_data[7]
port 484 nsew signal input
rlabel metal3 s 59200 43120 60000 43240 6 dcache_mem_o_data[8]
port 485 nsew signal input
rlabel metal3 s 59200 45568 60000 45688 6 dcache_mem_o_data[9]
port 486 nsew signal input
rlabel metal3 s 59200 17416 60000 17536 6 dcache_mem_req
port 487 nsew signal output
rlabel metal3 s 59200 22312 60000 22432 6 dcache_mem_sel[0]
port 488 nsew signal output
rlabel metal3 s 59200 25576 60000 25696 6 dcache_mem_sel[1]
port 489 nsew signal output
rlabel metal3 s 59200 17824 60000 17944 6 dcache_mem_we
port 490 nsew signal output
rlabel metal3 s 59200 18232 60000 18352 6 dcache_rst
port 491 nsew signal output
rlabel metal3 s 59200 18640 60000 18760 6 dcache_wb_4_burst
port 492 nsew signal input
rlabel metal3 s 59200 19048 60000 19168 6 dcache_wb_ack
port 493 nsew signal output
rlabel metal3 s 59200 22720 60000 22840 6 dcache_wb_adr[0]
port 494 nsew signal input
rlabel metal3 s 59200 48424 60000 48544 6 dcache_wb_adr[10]
port 495 nsew signal input
rlabel metal3 s 59200 50872 60000 50992 6 dcache_wb_adr[11]
port 496 nsew signal input
rlabel metal3 s 59200 53320 60000 53440 6 dcache_wb_adr[12]
port 497 nsew signal input
rlabel metal3 s 59200 55768 60000 55888 6 dcache_wb_adr[13]
port 498 nsew signal input
rlabel metal3 s 59200 58216 60000 58336 6 dcache_wb_adr[14]
port 499 nsew signal input
rlabel metal3 s 59200 60664 60000 60784 6 dcache_wb_adr[15]
port 500 nsew signal input
rlabel metal3 s 59200 62296 60000 62416 6 dcache_wb_adr[16]
port 501 nsew signal input
rlabel metal3 s 59200 63112 60000 63232 6 dcache_wb_adr[17]
port 502 nsew signal input
rlabel metal3 s 59200 63928 60000 64048 6 dcache_wb_adr[18]
port 503 nsew signal input
rlabel metal3 s 59200 64744 60000 64864 6 dcache_wb_adr[19]
port 504 nsew signal input
rlabel metal3 s 59200 25984 60000 26104 6 dcache_wb_adr[1]
port 505 nsew signal input
rlabel metal3 s 59200 65560 60000 65680 6 dcache_wb_adr[20]
port 506 nsew signal input
rlabel metal3 s 59200 66376 60000 66496 6 dcache_wb_adr[21]
port 507 nsew signal input
rlabel metal3 s 59200 67192 60000 67312 6 dcache_wb_adr[22]
port 508 nsew signal input
rlabel metal3 s 59200 68008 60000 68128 6 dcache_wb_adr[23]
port 509 nsew signal input
rlabel metal3 s 59200 28840 60000 28960 6 dcache_wb_adr[2]
port 510 nsew signal input
rlabel metal3 s 59200 31288 60000 31408 6 dcache_wb_adr[3]
port 511 nsew signal input
rlabel metal3 s 59200 33736 60000 33856 6 dcache_wb_adr[4]
port 512 nsew signal input
rlabel metal3 s 59200 36184 60000 36304 6 dcache_wb_adr[5]
port 513 nsew signal input
rlabel metal3 s 59200 38632 60000 38752 6 dcache_wb_adr[6]
port 514 nsew signal input
rlabel metal3 s 59200 41080 60000 41200 6 dcache_wb_adr[7]
port 515 nsew signal input
rlabel metal3 s 59200 43528 60000 43648 6 dcache_wb_adr[8]
port 516 nsew signal input
rlabel metal3 s 59200 45976 60000 46096 6 dcache_wb_adr[9]
port 517 nsew signal input
rlabel metal3 s 59200 19456 60000 19576 6 dcache_wb_cyc
port 518 nsew signal input
rlabel metal3 s 59200 19864 60000 19984 6 dcache_wb_err
port 519 nsew signal output
rlabel metal3 s 59200 23128 60000 23248 6 dcache_wb_i_dat[0]
port 520 nsew signal output
rlabel metal3 s 59200 48832 60000 48952 6 dcache_wb_i_dat[10]
port 521 nsew signal output
rlabel metal3 s 59200 51280 60000 51400 6 dcache_wb_i_dat[11]
port 522 nsew signal output
rlabel metal3 s 59200 53728 60000 53848 6 dcache_wb_i_dat[12]
port 523 nsew signal output
rlabel metal3 s 59200 56176 60000 56296 6 dcache_wb_i_dat[13]
port 524 nsew signal output
rlabel metal3 s 59200 58624 60000 58744 6 dcache_wb_i_dat[14]
port 525 nsew signal output
rlabel metal3 s 59200 61072 60000 61192 6 dcache_wb_i_dat[15]
port 526 nsew signal output
rlabel metal3 s 59200 26392 60000 26512 6 dcache_wb_i_dat[1]
port 527 nsew signal output
rlabel metal3 s 59200 29248 60000 29368 6 dcache_wb_i_dat[2]
port 528 nsew signal output
rlabel metal3 s 59200 31696 60000 31816 6 dcache_wb_i_dat[3]
port 529 nsew signal output
rlabel metal3 s 59200 34144 60000 34264 6 dcache_wb_i_dat[4]
port 530 nsew signal output
rlabel metal3 s 59200 36592 60000 36712 6 dcache_wb_i_dat[5]
port 531 nsew signal output
rlabel metal3 s 59200 39040 60000 39160 6 dcache_wb_i_dat[6]
port 532 nsew signal output
rlabel metal3 s 59200 41488 60000 41608 6 dcache_wb_i_dat[7]
port 533 nsew signal output
rlabel metal3 s 59200 43936 60000 44056 6 dcache_wb_i_dat[8]
port 534 nsew signal output
rlabel metal3 s 59200 46384 60000 46504 6 dcache_wb_i_dat[9]
port 535 nsew signal output
rlabel metal3 s 59200 23536 60000 23656 6 dcache_wb_o_dat[0]
port 536 nsew signal input
rlabel metal3 s 59200 49240 60000 49360 6 dcache_wb_o_dat[10]
port 537 nsew signal input
rlabel metal3 s 59200 51688 60000 51808 6 dcache_wb_o_dat[11]
port 538 nsew signal input
rlabel metal3 s 59200 54136 60000 54256 6 dcache_wb_o_dat[12]
port 539 nsew signal input
rlabel metal3 s 59200 56584 60000 56704 6 dcache_wb_o_dat[13]
port 540 nsew signal input
rlabel metal3 s 59200 59032 60000 59152 6 dcache_wb_o_dat[14]
port 541 nsew signal input
rlabel metal3 s 59200 61480 60000 61600 6 dcache_wb_o_dat[15]
port 542 nsew signal input
rlabel metal3 s 59200 26800 60000 26920 6 dcache_wb_o_dat[1]
port 543 nsew signal input
rlabel metal3 s 59200 29656 60000 29776 6 dcache_wb_o_dat[2]
port 544 nsew signal input
rlabel metal3 s 59200 32104 60000 32224 6 dcache_wb_o_dat[3]
port 545 nsew signal input
rlabel metal3 s 59200 34552 60000 34672 6 dcache_wb_o_dat[4]
port 546 nsew signal input
rlabel metal3 s 59200 37000 60000 37120 6 dcache_wb_o_dat[5]
port 547 nsew signal input
rlabel metal3 s 59200 39448 60000 39568 6 dcache_wb_o_dat[6]
port 548 nsew signal input
rlabel metal3 s 59200 41896 60000 42016 6 dcache_wb_o_dat[7]
port 549 nsew signal input
rlabel metal3 s 59200 44344 60000 44464 6 dcache_wb_o_dat[8]
port 550 nsew signal input
rlabel metal3 s 59200 46792 60000 46912 6 dcache_wb_o_dat[9]
port 551 nsew signal input
rlabel metal3 s 59200 23944 60000 24064 6 dcache_wb_sel[0]
port 552 nsew signal input
rlabel metal3 s 59200 27208 60000 27328 6 dcache_wb_sel[1]
port 553 nsew signal input
rlabel metal3 s 59200 20272 60000 20392 6 dcache_wb_stb
port 554 nsew signal input
rlabel metal3 s 59200 20680 60000 20800 6 dcache_wb_we
port 555 nsew signal input
rlabel metal3 s 59200 68416 60000 68536 6 ic0_clk
port 556 nsew signal output
rlabel metal3 s 59200 68824 60000 68944 6 ic0_mem_ack
port 557 nsew signal input
rlabel metal3 s 59200 72904 60000 73024 6 ic0_mem_addr[0]
port 558 nsew signal output
rlabel metal3 s 59200 90040 60000 90160 6 ic0_mem_addr[10]
port 559 nsew signal output
rlabel metal3 s 59200 91672 60000 91792 6 ic0_mem_addr[11]
port 560 nsew signal output
rlabel metal3 s 59200 93304 60000 93424 6 ic0_mem_addr[12]
port 561 nsew signal output
rlabel metal3 s 59200 94936 60000 95056 6 ic0_mem_addr[13]
port 562 nsew signal output
rlabel metal3 s 59200 96568 60000 96688 6 ic0_mem_addr[14]
port 563 nsew signal output
rlabel metal3 s 59200 98200 60000 98320 6 ic0_mem_addr[15]
port 564 nsew signal output
rlabel metal3 s 59200 74944 60000 75064 6 ic0_mem_addr[1]
port 565 nsew signal output
rlabel metal3 s 59200 76984 60000 77104 6 ic0_mem_addr[2]
port 566 nsew signal output
rlabel metal3 s 59200 78616 60000 78736 6 ic0_mem_addr[3]
port 567 nsew signal output
rlabel metal3 s 59200 80248 60000 80368 6 ic0_mem_addr[4]
port 568 nsew signal output
rlabel metal3 s 59200 81880 60000 82000 6 ic0_mem_addr[5]
port 569 nsew signal output
rlabel metal3 s 59200 83512 60000 83632 6 ic0_mem_addr[6]
port 570 nsew signal output
rlabel metal3 s 59200 85144 60000 85264 6 ic0_mem_addr[7]
port 571 nsew signal output
rlabel metal3 s 59200 86776 60000 86896 6 ic0_mem_addr[8]
port 572 nsew signal output
rlabel metal3 s 59200 88408 60000 88528 6 ic0_mem_addr[9]
port 573 nsew signal output
rlabel metal3 s 59200 69232 60000 69352 6 ic0_mem_cache_flush
port 574 nsew signal output
rlabel metal3 s 59200 73312 60000 73432 6 ic0_mem_data[0]
port 575 nsew signal input
rlabel metal3 s 59200 90448 60000 90568 6 ic0_mem_data[10]
port 576 nsew signal input
rlabel metal3 s 59200 92080 60000 92200 6 ic0_mem_data[11]
port 577 nsew signal input
rlabel metal3 s 59200 93712 60000 93832 6 ic0_mem_data[12]
port 578 nsew signal input
rlabel metal3 s 59200 95344 60000 95464 6 ic0_mem_data[13]
port 579 nsew signal input
rlabel metal3 s 59200 96976 60000 97096 6 ic0_mem_data[14]
port 580 nsew signal input
rlabel metal3 s 59200 98608 60000 98728 6 ic0_mem_data[15]
port 581 nsew signal input
rlabel metal3 s 59200 99832 60000 99952 6 ic0_mem_data[16]
port 582 nsew signal input
rlabel metal3 s 59200 100240 60000 100360 6 ic0_mem_data[17]
port 583 nsew signal input
rlabel metal3 s 59200 100648 60000 100768 6 ic0_mem_data[18]
port 584 nsew signal input
rlabel metal3 s 59200 101056 60000 101176 6 ic0_mem_data[19]
port 585 nsew signal input
rlabel metal3 s 59200 75352 60000 75472 6 ic0_mem_data[1]
port 586 nsew signal input
rlabel metal3 s 59200 101464 60000 101584 6 ic0_mem_data[20]
port 587 nsew signal input
rlabel metal3 s 59200 101872 60000 101992 6 ic0_mem_data[21]
port 588 nsew signal input
rlabel metal3 s 59200 102280 60000 102400 6 ic0_mem_data[22]
port 589 nsew signal input
rlabel metal3 s 59200 102688 60000 102808 6 ic0_mem_data[23]
port 590 nsew signal input
rlabel metal3 s 59200 103096 60000 103216 6 ic0_mem_data[24]
port 591 nsew signal input
rlabel metal3 s 59200 103504 60000 103624 6 ic0_mem_data[25]
port 592 nsew signal input
rlabel metal3 s 59200 103912 60000 104032 6 ic0_mem_data[26]
port 593 nsew signal input
rlabel metal3 s 59200 104320 60000 104440 6 ic0_mem_data[27]
port 594 nsew signal input
rlabel metal3 s 59200 104728 60000 104848 6 ic0_mem_data[28]
port 595 nsew signal input
rlabel metal3 s 59200 105136 60000 105256 6 ic0_mem_data[29]
port 596 nsew signal input
rlabel metal3 s 59200 77392 60000 77512 6 ic0_mem_data[2]
port 597 nsew signal input
rlabel metal3 s 59200 105544 60000 105664 6 ic0_mem_data[30]
port 598 nsew signal input
rlabel metal3 s 59200 105952 60000 106072 6 ic0_mem_data[31]
port 599 nsew signal input
rlabel metal3 s 59200 79024 60000 79144 6 ic0_mem_data[3]
port 600 nsew signal input
rlabel metal3 s 59200 80656 60000 80776 6 ic0_mem_data[4]
port 601 nsew signal input
rlabel metal3 s 59200 82288 60000 82408 6 ic0_mem_data[5]
port 602 nsew signal input
rlabel metal3 s 59200 83920 60000 84040 6 ic0_mem_data[6]
port 603 nsew signal input
rlabel metal3 s 59200 85552 60000 85672 6 ic0_mem_data[7]
port 604 nsew signal input
rlabel metal3 s 59200 87184 60000 87304 6 ic0_mem_data[8]
port 605 nsew signal input
rlabel metal3 s 59200 88816 60000 88936 6 ic0_mem_data[9]
port 606 nsew signal input
rlabel metal3 s 59200 69640 60000 69760 6 ic0_mem_ppl_submit
port 607 nsew signal output
rlabel metal3 s 59200 70048 60000 70168 6 ic0_mem_req
port 608 nsew signal output
rlabel metal3 s 59200 70456 60000 70576 6 ic0_rst
port 609 nsew signal output
rlabel metal3 s 59200 70864 60000 70984 6 ic0_wb_ack
port 610 nsew signal output
rlabel metal3 s 59200 73720 60000 73840 6 ic0_wb_adr[0]
port 611 nsew signal input
rlabel metal3 s 59200 90856 60000 90976 6 ic0_wb_adr[10]
port 612 nsew signal input
rlabel metal3 s 59200 92488 60000 92608 6 ic0_wb_adr[11]
port 613 nsew signal input
rlabel metal3 s 59200 94120 60000 94240 6 ic0_wb_adr[12]
port 614 nsew signal input
rlabel metal3 s 59200 95752 60000 95872 6 ic0_wb_adr[13]
port 615 nsew signal input
rlabel metal3 s 59200 97384 60000 97504 6 ic0_wb_adr[14]
port 616 nsew signal input
rlabel metal3 s 59200 99016 60000 99136 6 ic0_wb_adr[15]
port 617 nsew signal input
rlabel metal3 s 59200 75760 60000 75880 6 ic0_wb_adr[1]
port 618 nsew signal input
rlabel metal3 s 59200 77800 60000 77920 6 ic0_wb_adr[2]
port 619 nsew signal input
rlabel metal3 s 59200 79432 60000 79552 6 ic0_wb_adr[3]
port 620 nsew signal input
rlabel metal3 s 59200 81064 60000 81184 6 ic0_wb_adr[4]
port 621 nsew signal input
rlabel metal3 s 59200 82696 60000 82816 6 ic0_wb_adr[5]
port 622 nsew signal input
rlabel metal3 s 59200 84328 60000 84448 6 ic0_wb_adr[6]
port 623 nsew signal input
rlabel metal3 s 59200 85960 60000 86080 6 ic0_wb_adr[7]
port 624 nsew signal input
rlabel metal3 s 59200 87592 60000 87712 6 ic0_wb_adr[8]
port 625 nsew signal input
rlabel metal3 s 59200 89224 60000 89344 6 ic0_wb_adr[9]
port 626 nsew signal input
rlabel metal3 s 59200 71272 60000 71392 6 ic0_wb_cyc
port 627 nsew signal input
rlabel metal3 s 59200 71680 60000 71800 6 ic0_wb_err
port 628 nsew signal output
rlabel metal3 s 59200 74128 60000 74248 6 ic0_wb_i_dat[0]
port 629 nsew signal output
rlabel metal3 s 59200 91264 60000 91384 6 ic0_wb_i_dat[10]
port 630 nsew signal output
rlabel metal3 s 59200 92896 60000 93016 6 ic0_wb_i_dat[11]
port 631 nsew signal output
rlabel metal3 s 59200 94528 60000 94648 6 ic0_wb_i_dat[12]
port 632 nsew signal output
rlabel metal3 s 59200 96160 60000 96280 6 ic0_wb_i_dat[13]
port 633 nsew signal output
rlabel metal3 s 59200 97792 60000 97912 6 ic0_wb_i_dat[14]
port 634 nsew signal output
rlabel metal3 s 59200 99424 60000 99544 6 ic0_wb_i_dat[15]
port 635 nsew signal output
rlabel metal3 s 59200 76168 60000 76288 6 ic0_wb_i_dat[1]
port 636 nsew signal output
rlabel metal3 s 59200 78208 60000 78328 6 ic0_wb_i_dat[2]
port 637 nsew signal output
rlabel metal3 s 59200 79840 60000 79960 6 ic0_wb_i_dat[3]
port 638 nsew signal output
rlabel metal3 s 59200 81472 60000 81592 6 ic0_wb_i_dat[4]
port 639 nsew signal output
rlabel metal3 s 59200 83104 60000 83224 6 ic0_wb_i_dat[5]
port 640 nsew signal output
rlabel metal3 s 59200 84736 60000 84856 6 ic0_wb_i_dat[6]
port 641 nsew signal output
rlabel metal3 s 59200 86368 60000 86488 6 ic0_wb_i_dat[7]
port 642 nsew signal output
rlabel metal3 s 59200 88000 60000 88120 6 ic0_wb_i_dat[8]
port 643 nsew signal output
rlabel metal3 s 59200 89632 60000 89752 6 ic0_wb_i_dat[9]
port 644 nsew signal output
rlabel metal3 s 59200 74536 60000 74656 6 ic0_wb_sel[0]
port 645 nsew signal input
rlabel metal3 s 59200 76576 60000 76696 6 ic0_wb_sel[1]
port 646 nsew signal input
rlabel metal3 s 59200 72088 60000 72208 6 ic0_wb_stb
port 647 nsew signal input
rlabel metal3 s 59200 72496 60000 72616 6 ic0_wb_we
port 648 nsew signal input
rlabel metal3 s 59200 106360 60000 106480 6 ic1_clk
port 649 nsew signal output
rlabel metal3 s 59200 106768 60000 106888 6 ic1_mem_ack
port 650 nsew signal input
rlabel metal3 s 59200 110848 60000 110968 6 ic1_mem_addr[0]
port 651 nsew signal output
rlabel metal3 s 59200 127984 60000 128104 6 ic1_mem_addr[10]
port 652 nsew signal output
rlabel metal3 s 59200 129616 60000 129736 6 ic1_mem_addr[11]
port 653 nsew signal output
rlabel metal3 s 59200 131248 60000 131368 6 ic1_mem_addr[12]
port 654 nsew signal output
rlabel metal3 s 59200 132880 60000 133000 6 ic1_mem_addr[13]
port 655 nsew signal output
rlabel metal3 s 59200 134512 60000 134632 6 ic1_mem_addr[14]
port 656 nsew signal output
rlabel metal3 s 59200 136144 60000 136264 6 ic1_mem_addr[15]
port 657 nsew signal output
rlabel metal3 s 59200 112888 60000 113008 6 ic1_mem_addr[1]
port 658 nsew signal output
rlabel metal3 s 59200 114928 60000 115048 6 ic1_mem_addr[2]
port 659 nsew signal output
rlabel metal3 s 59200 116560 60000 116680 6 ic1_mem_addr[3]
port 660 nsew signal output
rlabel metal3 s 59200 118192 60000 118312 6 ic1_mem_addr[4]
port 661 nsew signal output
rlabel metal3 s 59200 119824 60000 119944 6 ic1_mem_addr[5]
port 662 nsew signal output
rlabel metal3 s 59200 121456 60000 121576 6 ic1_mem_addr[6]
port 663 nsew signal output
rlabel metal3 s 59200 123088 60000 123208 6 ic1_mem_addr[7]
port 664 nsew signal output
rlabel metal3 s 59200 124720 60000 124840 6 ic1_mem_addr[8]
port 665 nsew signal output
rlabel metal3 s 59200 126352 60000 126472 6 ic1_mem_addr[9]
port 666 nsew signal output
rlabel metal3 s 59200 107176 60000 107296 6 ic1_mem_cache_flush
port 667 nsew signal output
rlabel metal3 s 59200 111256 60000 111376 6 ic1_mem_data[0]
port 668 nsew signal input
rlabel metal3 s 59200 128392 60000 128512 6 ic1_mem_data[10]
port 669 nsew signal input
rlabel metal3 s 59200 130024 60000 130144 6 ic1_mem_data[11]
port 670 nsew signal input
rlabel metal3 s 59200 131656 60000 131776 6 ic1_mem_data[12]
port 671 nsew signal input
rlabel metal3 s 59200 133288 60000 133408 6 ic1_mem_data[13]
port 672 nsew signal input
rlabel metal3 s 59200 134920 60000 135040 6 ic1_mem_data[14]
port 673 nsew signal input
rlabel metal3 s 59200 136552 60000 136672 6 ic1_mem_data[15]
port 674 nsew signal input
rlabel metal3 s 59200 137776 60000 137896 6 ic1_mem_data[16]
port 675 nsew signal input
rlabel metal3 s 59200 138184 60000 138304 6 ic1_mem_data[17]
port 676 nsew signal input
rlabel metal3 s 59200 138592 60000 138712 6 ic1_mem_data[18]
port 677 nsew signal input
rlabel metal3 s 59200 139000 60000 139120 6 ic1_mem_data[19]
port 678 nsew signal input
rlabel metal3 s 59200 113296 60000 113416 6 ic1_mem_data[1]
port 679 nsew signal input
rlabel metal3 s 59200 139408 60000 139528 6 ic1_mem_data[20]
port 680 nsew signal input
rlabel metal3 s 59200 139816 60000 139936 6 ic1_mem_data[21]
port 681 nsew signal input
rlabel metal3 s 59200 140224 60000 140344 6 ic1_mem_data[22]
port 682 nsew signal input
rlabel metal3 s 59200 140632 60000 140752 6 ic1_mem_data[23]
port 683 nsew signal input
rlabel metal3 s 59200 141040 60000 141160 6 ic1_mem_data[24]
port 684 nsew signal input
rlabel metal3 s 59200 141448 60000 141568 6 ic1_mem_data[25]
port 685 nsew signal input
rlabel metal3 s 59200 141856 60000 141976 6 ic1_mem_data[26]
port 686 nsew signal input
rlabel metal3 s 59200 142264 60000 142384 6 ic1_mem_data[27]
port 687 nsew signal input
rlabel metal3 s 59200 142672 60000 142792 6 ic1_mem_data[28]
port 688 nsew signal input
rlabel metal3 s 59200 143080 60000 143200 6 ic1_mem_data[29]
port 689 nsew signal input
rlabel metal3 s 59200 115336 60000 115456 6 ic1_mem_data[2]
port 690 nsew signal input
rlabel metal3 s 59200 143488 60000 143608 6 ic1_mem_data[30]
port 691 nsew signal input
rlabel metal3 s 59200 143896 60000 144016 6 ic1_mem_data[31]
port 692 nsew signal input
rlabel metal3 s 59200 116968 60000 117088 6 ic1_mem_data[3]
port 693 nsew signal input
rlabel metal3 s 59200 118600 60000 118720 6 ic1_mem_data[4]
port 694 nsew signal input
rlabel metal3 s 59200 120232 60000 120352 6 ic1_mem_data[5]
port 695 nsew signal input
rlabel metal3 s 59200 121864 60000 121984 6 ic1_mem_data[6]
port 696 nsew signal input
rlabel metal3 s 59200 123496 60000 123616 6 ic1_mem_data[7]
port 697 nsew signal input
rlabel metal3 s 59200 125128 60000 125248 6 ic1_mem_data[8]
port 698 nsew signal input
rlabel metal3 s 59200 126760 60000 126880 6 ic1_mem_data[9]
port 699 nsew signal input
rlabel metal3 s 59200 107584 60000 107704 6 ic1_mem_ppl_submit
port 700 nsew signal output
rlabel metal3 s 59200 107992 60000 108112 6 ic1_mem_req
port 701 nsew signal output
rlabel metal3 s 59200 108400 60000 108520 6 ic1_rst
port 702 nsew signal output
rlabel metal3 s 59200 108808 60000 108928 6 ic1_wb_ack
port 703 nsew signal output
rlabel metal3 s 59200 111664 60000 111784 6 ic1_wb_adr[0]
port 704 nsew signal input
rlabel metal3 s 59200 128800 60000 128920 6 ic1_wb_adr[10]
port 705 nsew signal input
rlabel metal3 s 59200 130432 60000 130552 6 ic1_wb_adr[11]
port 706 nsew signal input
rlabel metal3 s 59200 132064 60000 132184 6 ic1_wb_adr[12]
port 707 nsew signal input
rlabel metal3 s 59200 133696 60000 133816 6 ic1_wb_adr[13]
port 708 nsew signal input
rlabel metal3 s 59200 135328 60000 135448 6 ic1_wb_adr[14]
port 709 nsew signal input
rlabel metal3 s 59200 136960 60000 137080 6 ic1_wb_adr[15]
port 710 nsew signal input
rlabel metal3 s 59200 113704 60000 113824 6 ic1_wb_adr[1]
port 711 nsew signal input
rlabel metal3 s 59200 115744 60000 115864 6 ic1_wb_adr[2]
port 712 nsew signal input
rlabel metal3 s 59200 117376 60000 117496 6 ic1_wb_adr[3]
port 713 nsew signal input
rlabel metal3 s 59200 119008 60000 119128 6 ic1_wb_adr[4]
port 714 nsew signal input
rlabel metal3 s 59200 120640 60000 120760 6 ic1_wb_adr[5]
port 715 nsew signal input
rlabel metal3 s 59200 122272 60000 122392 6 ic1_wb_adr[6]
port 716 nsew signal input
rlabel metal3 s 59200 123904 60000 124024 6 ic1_wb_adr[7]
port 717 nsew signal input
rlabel metal3 s 59200 125536 60000 125656 6 ic1_wb_adr[8]
port 718 nsew signal input
rlabel metal3 s 59200 127168 60000 127288 6 ic1_wb_adr[9]
port 719 nsew signal input
rlabel metal3 s 59200 109216 60000 109336 6 ic1_wb_cyc
port 720 nsew signal input
rlabel metal3 s 59200 109624 60000 109744 6 ic1_wb_err
port 721 nsew signal output
rlabel metal3 s 59200 112072 60000 112192 6 ic1_wb_i_dat[0]
port 722 nsew signal output
rlabel metal3 s 59200 129208 60000 129328 6 ic1_wb_i_dat[10]
port 723 nsew signal output
rlabel metal3 s 59200 130840 60000 130960 6 ic1_wb_i_dat[11]
port 724 nsew signal output
rlabel metal3 s 59200 132472 60000 132592 6 ic1_wb_i_dat[12]
port 725 nsew signal output
rlabel metal3 s 59200 134104 60000 134224 6 ic1_wb_i_dat[13]
port 726 nsew signal output
rlabel metal3 s 59200 135736 60000 135856 6 ic1_wb_i_dat[14]
port 727 nsew signal output
rlabel metal3 s 59200 137368 60000 137488 6 ic1_wb_i_dat[15]
port 728 nsew signal output
rlabel metal3 s 59200 114112 60000 114232 6 ic1_wb_i_dat[1]
port 729 nsew signal output
rlabel metal3 s 59200 116152 60000 116272 6 ic1_wb_i_dat[2]
port 730 nsew signal output
rlabel metal3 s 59200 117784 60000 117904 6 ic1_wb_i_dat[3]
port 731 nsew signal output
rlabel metal3 s 59200 119416 60000 119536 6 ic1_wb_i_dat[4]
port 732 nsew signal output
rlabel metal3 s 59200 121048 60000 121168 6 ic1_wb_i_dat[5]
port 733 nsew signal output
rlabel metal3 s 59200 122680 60000 122800 6 ic1_wb_i_dat[6]
port 734 nsew signal output
rlabel metal3 s 59200 124312 60000 124432 6 ic1_wb_i_dat[7]
port 735 nsew signal output
rlabel metal3 s 59200 125944 60000 126064 6 ic1_wb_i_dat[8]
port 736 nsew signal output
rlabel metal3 s 59200 127576 60000 127696 6 ic1_wb_i_dat[9]
port 737 nsew signal output
rlabel metal3 s 59200 112480 60000 112600 6 ic1_wb_sel[0]
port 738 nsew signal input
rlabel metal3 s 59200 114520 60000 114640 6 ic1_wb_sel[1]
port 739 nsew signal input
rlabel metal3 s 59200 110032 60000 110152 6 ic1_wb_stb
port 740 nsew signal input
rlabel metal3 s 59200 110440 60000 110560 6 ic1_wb_we
port 741 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 inner_disable
port 742 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 inner_embed_mode
port 743 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 inner_ext_irq
port 744 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 inner_wb_4_burst
port 745 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 inner_wb_8_burst
port 746 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 inner_wb_ack
port 747 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 inner_wb_adr[0]
port 748 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 inner_wb_adr[10]
port 749 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 inner_wb_adr[11]
port 750 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 inner_wb_adr[12]
port 751 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 inner_wb_adr[13]
port 752 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 inner_wb_adr[14]
port 753 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 inner_wb_adr[15]
port 754 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 inner_wb_adr[16]
port 755 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 inner_wb_adr[17]
port 756 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 inner_wb_adr[18]
port 757 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 inner_wb_adr[19]
port 758 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 inner_wb_adr[1]
port 759 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 inner_wb_adr[20]
port 760 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 inner_wb_adr[21]
port 761 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 inner_wb_adr[22]
port 762 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 inner_wb_adr[23]
port 763 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 inner_wb_adr[2]
port 764 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 inner_wb_adr[3]
port 765 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 inner_wb_adr[4]
port 766 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 inner_wb_adr[5]
port 767 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 inner_wb_adr[6]
port 768 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 inner_wb_adr[7]
port 769 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 inner_wb_adr[8]
port 770 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 inner_wb_adr[9]
port 771 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 inner_wb_cyc
port 772 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 inner_wb_err
port 773 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 inner_wb_i_dat[0]
port 774 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 inner_wb_i_dat[10]
port 775 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 inner_wb_i_dat[11]
port 776 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 inner_wb_i_dat[12]
port 777 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 inner_wb_i_dat[13]
port 778 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 inner_wb_i_dat[14]
port 779 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 inner_wb_i_dat[15]
port 780 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 inner_wb_i_dat[1]
port 781 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 inner_wb_i_dat[2]
port 782 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 inner_wb_i_dat[3]
port 783 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 inner_wb_i_dat[4]
port 784 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 inner_wb_i_dat[5]
port 785 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 inner_wb_i_dat[6]
port 786 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 inner_wb_i_dat[7]
port 787 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 inner_wb_i_dat[8]
port 788 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 inner_wb_i_dat[9]
port 789 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 inner_wb_o_dat[0]
port 790 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 inner_wb_o_dat[10]
port 791 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 inner_wb_o_dat[11]
port 792 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 inner_wb_o_dat[12]
port 793 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 inner_wb_o_dat[13]
port 794 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 inner_wb_o_dat[14]
port 795 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 inner_wb_o_dat[15]
port 796 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 inner_wb_o_dat[1]
port 797 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 inner_wb_o_dat[2]
port 798 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 inner_wb_o_dat[3]
port 799 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 inner_wb_o_dat[4]
port 800 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 inner_wb_o_dat[5]
port 801 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 inner_wb_o_dat[6]
port 802 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 inner_wb_o_dat[7]
port 803 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 inner_wb_o_dat[8]
port 804 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 inner_wb_o_dat[9]
port 805 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 inner_wb_sel[0]
port 806 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 inner_wb_sel[1]
port 807 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 inner_wb_stb
port 808 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 inner_wb_we
port 809 nsew signal output
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 810 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 810 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 811 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 811 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 20219510
string GDS_FILE /home/piotro/caravel_user_project/openlane/interconnect_inner/runs/22_12_30_18_27/results/signoff/interconnect_inner.magic.gds
string GDS_START 857996
<< end >>

