magic
tech gf180mcuD
magscale 1 5
timestamp 1699782230
<< obsm1 >>
rect 672 1538 49280 98881
<< metal2 >>
rect 1344 99600 1400 100000
rect 1568 99600 1624 100000
rect 1792 99600 1848 100000
rect 2016 99600 2072 100000
rect 2240 99600 2296 100000
rect 2464 99600 2520 100000
rect 2688 99600 2744 100000
rect 2912 99600 2968 100000
rect 3136 99600 3192 100000
rect 3360 99600 3416 100000
rect 3584 99600 3640 100000
rect 3808 99600 3864 100000
rect 4032 99600 4088 100000
rect 4256 99600 4312 100000
rect 4480 99600 4536 100000
rect 4704 99600 4760 100000
rect 4928 99600 4984 100000
rect 5152 99600 5208 100000
rect 5376 99600 5432 100000
rect 5600 99600 5656 100000
rect 5824 99600 5880 100000
rect 6048 99600 6104 100000
rect 6272 99600 6328 100000
rect 6496 99600 6552 100000
rect 6720 99600 6776 100000
rect 6944 99600 7000 100000
rect 7168 99600 7224 100000
rect 7392 99600 7448 100000
rect 7616 99600 7672 100000
rect 7840 99600 7896 100000
rect 8064 99600 8120 100000
rect 8288 99600 8344 100000
rect 8512 99600 8568 100000
rect 8736 99600 8792 100000
rect 8960 99600 9016 100000
rect 9184 99600 9240 100000
rect 9408 99600 9464 100000
rect 9632 99600 9688 100000
rect 9856 99600 9912 100000
rect 10080 99600 10136 100000
rect 10304 99600 10360 100000
rect 10528 99600 10584 100000
rect 10752 99600 10808 100000
rect 10976 99600 11032 100000
rect 11200 99600 11256 100000
rect 11424 99600 11480 100000
rect 11648 99600 11704 100000
rect 11872 99600 11928 100000
rect 12096 99600 12152 100000
rect 12320 99600 12376 100000
rect 12544 99600 12600 100000
rect 12768 99600 12824 100000
rect 12992 99600 13048 100000
rect 13216 99600 13272 100000
rect 13440 99600 13496 100000
rect 13664 99600 13720 100000
rect 13888 99600 13944 100000
rect 14112 99600 14168 100000
rect 14336 99600 14392 100000
rect 14560 99600 14616 100000
rect 14784 99600 14840 100000
rect 15008 99600 15064 100000
rect 15232 99600 15288 100000
rect 15456 99600 15512 100000
rect 15680 99600 15736 100000
rect 15904 99600 15960 100000
rect 16128 99600 16184 100000
rect 16352 99600 16408 100000
rect 16576 99600 16632 100000
rect 16800 99600 16856 100000
rect 17024 99600 17080 100000
rect 17248 99600 17304 100000
rect 17472 99600 17528 100000
rect 17696 99600 17752 100000
rect 17920 99600 17976 100000
rect 18144 99600 18200 100000
rect 18368 99600 18424 100000
rect 18592 99600 18648 100000
rect 18816 99600 18872 100000
rect 19040 99600 19096 100000
rect 19264 99600 19320 100000
rect 19488 99600 19544 100000
rect 19712 99600 19768 100000
rect 19936 99600 19992 100000
rect 20160 99600 20216 100000
rect 20384 99600 20440 100000
rect 20608 99600 20664 100000
rect 20832 99600 20888 100000
rect 21056 99600 21112 100000
rect 21280 99600 21336 100000
rect 21504 99600 21560 100000
rect 21728 99600 21784 100000
rect 21952 99600 22008 100000
rect 22176 99600 22232 100000
rect 22400 99600 22456 100000
rect 22624 99600 22680 100000
rect 22848 99600 22904 100000
rect 23072 99600 23128 100000
rect 23296 99600 23352 100000
rect 23520 99600 23576 100000
rect 23744 99600 23800 100000
rect 23968 99600 24024 100000
rect 24192 99600 24248 100000
rect 24416 99600 24472 100000
rect 24640 99600 24696 100000
rect 24864 99600 24920 100000
rect 25088 99600 25144 100000
rect 25312 99600 25368 100000
rect 25536 99600 25592 100000
rect 25760 99600 25816 100000
rect 25984 99600 26040 100000
rect 26208 99600 26264 100000
rect 26432 99600 26488 100000
rect 26656 99600 26712 100000
rect 26880 99600 26936 100000
rect 27104 99600 27160 100000
rect 27328 99600 27384 100000
rect 27552 99600 27608 100000
rect 27776 99600 27832 100000
rect 28000 99600 28056 100000
rect 28224 99600 28280 100000
rect 28448 99600 28504 100000
rect 28672 99600 28728 100000
rect 28896 99600 28952 100000
rect 29120 99600 29176 100000
rect 29344 99600 29400 100000
rect 29568 99600 29624 100000
rect 29792 99600 29848 100000
rect 30016 99600 30072 100000
rect 30240 99600 30296 100000
rect 30464 99600 30520 100000
rect 30688 99600 30744 100000
rect 30912 99600 30968 100000
rect 31136 99600 31192 100000
rect 31360 99600 31416 100000
rect 31584 99600 31640 100000
rect 31808 99600 31864 100000
rect 32032 99600 32088 100000
rect 32256 99600 32312 100000
rect 32480 99600 32536 100000
rect 32704 99600 32760 100000
rect 32928 99600 32984 100000
rect 33152 99600 33208 100000
rect 33376 99600 33432 100000
rect 33600 99600 33656 100000
rect 33824 99600 33880 100000
rect 34048 99600 34104 100000
rect 34272 99600 34328 100000
rect 34496 99600 34552 100000
rect 34720 99600 34776 100000
rect 34944 99600 35000 100000
rect 35168 99600 35224 100000
rect 35392 99600 35448 100000
rect 35616 99600 35672 100000
rect 35840 99600 35896 100000
rect 36064 99600 36120 100000
rect 36288 99600 36344 100000
rect 36512 99600 36568 100000
rect 36736 99600 36792 100000
rect 36960 99600 37016 100000
rect 37184 99600 37240 100000
rect 37408 99600 37464 100000
rect 37632 99600 37688 100000
rect 37856 99600 37912 100000
rect 38080 99600 38136 100000
rect 38304 99600 38360 100000
rect 38528 99600 38584 100000
rect 38752 99600 38808 100000
rect 38976 99600 39032 100000
rect 39200 99600 39256 100000
rect 39424 99600 39480 100000
rect 39648 99600 39704 100000
rect 39872 99600 39928 100000
rect 40096 99600 40152 100000
rect 40320 99600 40376 100000
rect 40544 99600 40600 100000
rect 40768 99600 40824 100000
rect 40992 99600 41048 100000
rect 41216 99600 41272 100000
rect 41440 99600 41496 100000
rect 41664 99600 41720 100000
rect 41888 99600 41944 100000
rect 42112 99600 42168 100000
rect 42336 99600 42392 100000
rect 42560 99600 42616 100000
rect 42784 99600 42840 100000
rect 43008 99600 43064 100000
rect 43232 99600 43288 100000
rect 43456 99600 43512 100000
rect 43680 99600 43736 100000
rect 43904 99600 43960 100000
rect 44128 99600 44184 100000
rect 44352 99600 44408 100000
rect 44576 99600 44632 100000
rect 44800 99600 44856 100000
rect 45024 99600 45080 100000
rect 45248 99600 45304 100000
rect 45472 99600 45528 100000
rect 45696 99600 45752 100000
rect 45920 99600 45976 100000
rect 46144 99600 46200 100000
rect 46368 99600 46424 100000
rect 46592 99600 46648 100000
rect 46816 99600 46872 100000
rect 47040 99600 47096 100000
rect 47264 99600 47320 100000
rect 47488 99600 47544 100000
rect 47712 99600 47768 100000
rect 47936 99600 47992 100000
rect 48160 99600 48216 100000
rect 48384 99600 48440 100000
rect 48608 99600 48664 100000
<< obsm2 >>
rect 518 99570 1314 99600
rect 1430 99570 1538 99600
rect 1654 99570 1762 99600
rect 1878 99570 1986 99600
rect 2102 99570 2210 99600
rect 2326 99570 2434 99600
rect 2550 99570 2658 99600
rect 2774 99570 2882 99600
rect 2998 99570 3106 99600
rect 3222 99570 3330 99600
rect 3446 99570 3554 99600
rect 3670 99570 3778 99600
rect 3894 99570 4002 99600
rect 4118 99570 4226 99600
rect 4342 99570 4450 99600
rect 4566 99570 4674 99600
rect 4790 99570 4898 99600
rect 5014 99570 5122 99600
rect 5238 99570 5346 99600
rect 5462 99570 5570 99600
rect 5686 99570 5794 99600
rect 5910 99570 6018 99600
rect 6134 99570 6242 99600
rect 6358 99570 6466 99600
rect 6582 99570 6690 99600
rect 6806 99570 6914 99600
rect 7030 99570 7138 99600
rect 7254 99570 7362 99600
rect 7478 99570 7586 99600
rect 7702 99570 7810 99600
rect 7926 99570 8034 99600
rect 8150 99570 8258 99600
rect 8374 99570 8482 99600
rect 8598 99570 8706 99600
rect 8822 99570 8930 99600
rect 9046 99570 9154 99600
rect 9270 99570 9378 99600
rect 9494 99570 9602 99600
rect 9718 99570 9826 99600
rect 9942 99570 10050 99600
rect 10166 99570 10274 99600
rect 10390 99570 10498 99600
rect 10614 99570 10722 99600
rect 10838 99570 10946 99600
rect 11062 99570 11170 99600
rect 11286 99570 11394 99600
rect 11510 99570 11618 99600
rect 11734 99570 11842 99600
rect 11958 99570 12066 99600
rect 12182 99570 12290 99600
rect 12406 99570 12514 99600
rect 12630 99570 12738 99600
rect 12854 99570 12962 99600
rect 13078 99570 13186 99600
rect 13302 99570 13410 99600
rect 13526 99570 13634 99600
rect 13750 99570 13858 99600
rect 13974 99570 14082 99600
rect 14198 99570 14306 99600
rect 14422 99570 14530 99600
rect 14646 99570 14754 99600
rect 14870 99570 14978 99600
rect 15094 99570 15202 99600
rect 15318 99570 15426 99600
rect 15542 99570 15650 99600
rect 15766 99570 15874 99600
rect 15990 99570 16098 99600
rect 16214 99570 16322 99600
rect 16438 99570 16546 99600
rect 16662 99570 16770 99600
rect 16886 99570 16994 99600
rect 17110 99570 17218 99600
rect 17334 99570 17442 99600
rect 17558 99570 17666 99600
rect 17782 99570 17890 99600
rect 18006 99570 18114 99600
rect 18230 99570 18338 99600
rect 18454 99570 18562 99600
rect 18678 99570 18786 99600
rect 18902 99570 19010 99600
rect 19126 99570 19234 99600
rect 19350 99570 19458 99600
rect 19574 99570 19682 99600
rect 19798 99570 19906 99600
rect 20022 99570 20130 99600
rect 20246 99570 20354 99600
rect 20470 99570 20578 99600
rect 20694 99570 20802 99600
rect 20918 99570 21026 99600
rect 21142 99570 21250 99600
rect 21366 99570 21474 99600
rect 21590 99570 21698 99600
rect 21814 99570 21922 99600
rect 22038 99570 22146 99600
rect 22262 99570 22370 99600
rect 22486 99570 22594 99600
rect 22710 99570 22818 99600
rect 22934 99570 23042 99600
rect 23158 99570 23266 99600
rect 23382 99570 23490 99600
rect 23606 99570 23714 99600
rect 23830 99570 23938 99600
rect 24054 99570 24162 99600
rect 24278 99570 24386 99600
rect 24502 99570 24610 99600
rect 24726 99570 24834 99600
rect 24950 99570 25058 99600
rect 25174 99570 25282 99600
rect 25398 99570 25506 99600
rect 25622 99570 25730 99600
rect 25846 99570 25954 99600
rect 26070 99570 26178 99600
rect 26294 99570 26402 99600
rect 26518 99570 26626 99600
rect 26742 99570 26850 99600
rect 26966 99570 27074 99600
rect 27190 99570 27298 99600
rect 27414 99570 27522 99600
rect 27638 99570 27746 99600
rect 27862 99570 27970 99600
rect 28086 99570 28194 99600
rect 28310 99570 28418 99600
rect 28534 99570 28642 99600
rect 28758 99570 28866 99600
rect 28982 99570 29090 99600
rect 29206 99570 29314 99600
rect 29430 99570 29538 99600
rect 29654 99570 29762 99600
rect 29878 99570 29986 99600
rect 30102 99570 30210 99600
rect 30326 99570 30434 99600
rect 30550 99570 30658 99600
rect 30774 99570 30882 99600
rect 30998 99570 31106 99600
rect 31222 99570 31330 99600
rect 31446 99570 31554 99600
rect 31670 99570 31778 99600
rect 31894 99570 32002 99600
rect 32118 99570 32226 99600
rect 32342 99570 32450 99600
rect 32566 99570 32674 99600
rect 32790 99570 32898 99600
rect 33014 99570 33122 99600
rect 33238 99570 33346 99600
rect 33462 99570 33570 99600
rect 33686 99570 33794 99600
rect 33910 99570 34018 99600
rect 34134 99570 34242 99600
rect 34358 99570 34466 99600
rect 34582 99570 34690 99600
rect 34806 99570 34914 99600
rect 35030 99570 35138 99600
rect 35254 99570 35362 99600
rect 35478 99570 35586 99600
rect 35702 99570 35810 99600
rect 35926 99570 36034 99600
rect 36150 99570 36258 99600
rect 36374 99570 36482 99600
rect 36598 99570 36706 99600
rect 36822 99570 36930 99600
rect 37046 99570 37154 99600
rect 37270 99570 37378 99600
rect 37494 99570 37602 99600
rect 37718 99570 37826 99600
rect 37942 99570 38050 99600
rect 38166 99570 38274 99600
rect 38390 99570 38498 99600
rect 38614 99570 38722 99600
rect 38838 99570 38946 99600
rect 39062 99570 39170 99600
rect 39286 99570 39394 99600
rect 39510 99570 39618 99600
rect 39734 99570 39842 99600
rect 39958 99570 40066 99600
rect 40182 99570 40290 99600
rect 40406 99570 40514 99600
rect 40630 99570 40738 99600
rect 40854 99570 40962 99600
rect 41078 99570 41186 99600
rect 41302 99570 41410 99600
rect 41526 99570 41634 99600
rect 41750 99570 41858 99600
rect 41974 99570 42082 99600
rect 42198 99570 42306 99600
rect 42422 99570 42530 99600
rect 42646 99570 42754 99600
rect 42870 99570 42978 99600
rect 43094 99570 43202 99600
rect 43318 99570 43426 99600
rect 43542 99570 43650 99600
rect 43766 99570 43874 99600
rect 43990 99570 44098 99600
rect 44214 99570 44322 99600
rect 44438 99570 44546 99600
rect 44662 99570 44770 99600
rect 44886 99570 44994 99600
rect 45110 99570 45218 99600
rect 45334 99570 45442 99600
rect 45558 99570 45666 99600
rect 45782 99570 45890 99600
rect 46006 99570 46114 99600
rect 46230 99570 46338 99600
rect 46454 99570 46562 99600
rect 46678 99570 46786 99600
rect 46902 99570 47010 99600
rect 47126 99570 47234 99600
rect 47350 99570 47458 99600
rect 47574 99570 47682 99600
rect 47798 99570 47906 99600
rect 48022 99570 48130 99600
rect 48246 99570 48354 99600
rect 48470 99570 48578 99600
rect 48694 99570 49154 99600
rect 518 1549 49154 99570
<< obsm3 >>
rect 513 1554 49159 98602
<< metal4 >>
rect 2224 1538 2384 98422
rect 9904 1538 10064 98422
rect 17584 1538 17744 98422
rect 25264 1538 25424 98422
rect 32944 1538 33104 98422
rect 40624 1538 40784 98422
rect 48304 1538 48464 98422
<< obsm4 >>
rect 2702 3033 9874 98103
rect 10094 3033 17554 98103
rect 17774 3033 25234 98103
rect 25454 3033 32914 98103
rect 33134 3033 40594 98103
rect 40814 3033 47306 98103
<< labels >>
rlabel metal2 s 5376 99600 5432 100000 6 dbg_pc[0]
port 1 nsew signal output
rlabel metal2 s 31808 99600 31864 100000 6 dbg_pc[10]
port 2 nsew signal output
rlabel metal2 s 34048 99600 34104 100000 6 dbg_pc[11]
port 3 nsew signal output
rlabel metal2 s 36288 99600 36344 100000 6 dbg_pc[12]
port 4 nsew signal output
rlabel metal2 s 38528 99600 38584 100000 6 dbg_pc[13]
port 5 nsew signal output
rlabel metal2 s 40768 99600 40824 100000 6 dbg_pc[14]
port 6 nsew signal output
rlabel metal2 s 43008 99600 43064 100000 6 dbg_pc[15]
port 7 nsew signal output
rlabel metal2 s 8288 99600 8344 100000 6 dbg_pc[1]
port 8 nsew signal output
rlabel metal2 s 11200 99600 11256 100000 6 dbg_pc[2]
port 9 nsew signal output
rlabel metal2 s 13888 99600 13944 100000 6 dbg_pc[3]
port 10 nsew signal output
rlabel metal2 s 16576 99600 16632 100000 6 dbg_pc[4]
port 11 nsew signal output
rlabel metal2 s 19264 99600 19320 100000 6 dbg_pc[5]
port 12 nsew signal output
rlabel metal2 s 21952 99600 22008 100000 6 dbg_pc[6]
port 13 nsew signal output
rlabel metal2 s 24640 99600 24696 100000 6 dbg_pc[7]
port 14 nsew signal output
rlabel metal2 s 27328 99600 27384 100000 6 dbg_pc[8]
port 15 nsew signal output
rlabel metal2 s 29568 99600 29624 100000 6 dbg_pc[9]
port 16 nsew signal output
rlabel metal2 s 5600 99600 5656 100000 6 dbg_r0[0]
port 17 nsew signal output
rlabel metal2 s 32032 99600 32088 100000 6 dbg_r0[10]
port 18 nsew signal output
rlabel metal2 s 34272 99600 34328 100000 6 dbg_r0[11]
port 19 nsew signal output
rlabel metal2 s 36512 99600 36568 100000 6 dbg_r0[12]
port 20 nsew signal output
rlabel metal2 s 38752 99600 38808 100000 6 dbg_r0[13]
port 21 nsew signal output
rlabel metal2 s 40992 99600 41048 100000 6 dbg_r0[14]
port 22 nsew signal output
rlabel metal2 s 43232 99600 43288 100000 6 dbg_r0[15]
port 23 nsew signal output
rlabel metal2 s 8512 99600 8568 100000 6 dbg_r0[1]
port 24 nsew signal output
rlabel metal2 s 11424 99600 11480 100000 6 dbg_r0[2]
port 25 nsew signal output
rlabel metal2 s 14112 99600 14168 100000 6 dbg_r0[3]
port 26 nsew signal output
rlabel metal2 s 16800 99600 16856 100000 6 dbg_r0[4]
port 27 nsew signal output
rlabel metal2 s 19488 99600 19544 100000 6 dbg_r0[5]
port 28 nsew signal output
rlabel metal2 s 22176 99600 22232 100000 6 dbg_r0[6]
port 29 nsew signal output
rlabel metal2 s 24864 99600 24920 100000 6 dbg_r0[7]
port 30 nsew signal output
rlabel metal2 s 27552 99600 27608 100000 6 dbg_r0[8]
port 31 nsew signal output
rlabel metal2 s 29792 99600 29848 100000 6 dbg_r0[9]
port 32 nsew signal output
rlabel metal2 s 1344 99600 1400 100000 6 i_clk
port 33 nsew signal input
rlabel metal2 s 5824 99600 5880 100000 6 i_core_int_sreg[0]
port 34 nsew signal input
rlabel metal2 s 32256 99600 32312 100000 6 i_core_int_sreg[10]
port 35 nsew signal input
rlabel metal2 s 34496 99600 34552 100000 6 i_core_int_sreg[11]
port 36 nsew signal input
rlabel metal2 s 36736 99600 36792 100000 6 i_core_int_sreg[12]
port 37 nsew signal input
rlabel metal2 s 38976 99600 39032 100000 6 i_core_int_sreg[13]
port 38 nsew signal input
rlabel metal2 s 41216 99600 41272 100000 6 i_core_int_sreg[14]
port 39 nsew signal input
rlabel metal2 s 43456 99600 43512 100000 6 i_core_int_sreg[15]
port 40 nsew signal input
rlabel metal2 s 8736 99600 8792 100000 6 i_core_int_sreg[1]
port 41 nsew signal input
rlabel metal2 s 11648 99600 11704 100000 6 i_core_int_sreg[2]
port 42 nsew signal input
rlabel metal2 s 14336 99600 14392 100000 6 i_core_int_sreg[3]
port 43 nsew signal input
rlabel metal2 s 17024 99600 17080 100000 6 i_core_int_sreg[4]
port 44 nsew signal input
rlabel metal2 s 19712 99600 19768 100000 6 i_core_int_sreg[5]
port 45 nsew signal input
rlabel metal2 s 22400 99600 22456 100000 6 i_core_int_sreg[6]
port 46 nsew signal input
rlabel metal2 s 25088 99600 25144 100000 6 i_core_int_sreg[7]
port 47 nsew signal input
rlabel metal2 s 27776 99600 27832 100000 6 i_core_int_sreg[8]
port 48 nsew signal input
rlabel metal2 s 30016 99600 30072 100000 6 i_core_int_sreg[9]
port 49 nsew signal input
rlabel metal2 s 1568 99600 1624 100000 6 i_disable
port 50 nsew signal input
rlabel metal2 s 1792 99600 1848 100000 6 i_irq
port 51 nsew signal input
rlabel metal2 s 2016 99600 2072 100000 6 i_mc_core_int
port 52 nsew signal input
rlabel metal2 s 2240 99600 2296 100000 6 i_mem_ack
port 53 nsew signal input
rlabel metal2 s 6048 99600 6104 100000 6 i_mem_data[0]
port 54 nsew signal input
rlabel metal2 s 32480 99600 32536 100000 6 i_mem_data[10]
port 55 nsew signal input
rlabel metal2 s 34720 99600 34776 100000 6 i_mem_data[11]
port 56 nsew signal input
rlabel metal2 s 36960 99600 37016 100000 6 i_mem_data[12]
port 57 nsew signal input
rlabel metal2 s 39200 99600 39256 100000 6 i_mem_data[13]
port 58 nsew signal input
rlabel metal2 s 41440 99600 41496 100000 6 i_mem_data[14]
port 59 nsew signal input
rlabel metal2 s 43680 99600 43736 100000 6 i_mem_data[15]
port 60 nsew signal input
rlabel metal2 s 8960 99600 9016 100000 6 i_mem_data[1]
port 61 nsew signal input
rlabel metal2 s 11872 99600 11928 100000 6 i_mem_data[2]
port 62 nsew signal input
rlabel metal2 s 14560 99600 14616 100000 6 i_mem_data[3]
port 63 nsew signal input
rlabel metal2 s 17248 99600 17304 100000 6 i_mem_data[4]
port 64 nsew signal input
rlabel metal2 s 19936 99600 19992 100000 6 i_mem_data[5]
port 65 nsew signal input
rlabel metal2 s 22624 99600 22680 100000 6 i_mem_data[6]
port 66 nsew signal input
rlabel metal2 s 25312 99600 25368 100000 6 i_mem_data[7]
port 67 nsew signal input
rlabel metal2 s 28000 99600 28056 100000 6 i_mem_data[8]
port 68 nsew signal input
rlabel metal2 s 30240 99600 30296 100000 6 i_mem_data[9]
port 69 nsew signal input
rlabel metal2 s 2464 99600 2520 100000 6 i_mem_exception
port 70 nsew signal input
rlabel metal2 s 6272 99600 6328 100000 6 i_req_data[0]
port 71 nsew signal input
rlabel metal2 s 32704 99600 32760 100000 6 i_req_data[10]
port 72 nsew signal input
rlabel metal2 s 34944 99600 35000 100000 6 i_req_data[11]
port 73 nsew signal input
rlabel metal2 s 37184 99600 37240 100000 6 i_req_data[12]
port 74 nsew signal input
rlabel metal2 s 39424 99600 39480 100000 6 i_req_data[13]
port 75 nsew signal input
rlabel metal2 s 41664 99600 41720 100000 6 i_req_data[14]
port 76 nsew signal input
rlabel metal2 s 43904 99600 43960 100000 6 i_req_data[15]
port 77 nsew signal input
rlabel metal2 s 45248 99600 45304 100000 6 i_req_data[16]
port 78 nsew signal input
rlabel metal2 s 45472 99600 45528 100000 6 i_req_data[17]
port 79 nsew signal input
rlabel metal2 s 45696 99600 45752 100000 6 i_req_data[18]
port 80 nsew signal input
rlabel metal2 s 45920 99600 45976 100000 6 i_req_data[19]
port 81 nsew signal input
rlabel metal2 s 9184 99600 9240 100000 6 i_req_data[1]
port 82 nsew signal input
rlabel metal2 s 46144 99600 46200 100000 6 i_req_data[20]
port 83 nsew signal input
rlabel metal2 s 46368 99600 46424 100000 6 i_req_data[21]
port 84 nsew signal input
rlabel metal2 s 46592 99600 46648 100000 6 i_req_data[22]
port 85 nsew signal input
rlabel metal2 s 46816 99600 46872 100000 6 i_req_data[23]
port 86 nsew signal input
rlabel metal2 s 47040 99600 47096 100000 6 i_req_data[24]
port 87 nsew signal input
rlabel metal2 s 47264 99600 47320 100000 6 i_req_data[25]
port 88 nsew signal input
rlabel metal2 s 47488 99600 47544 100000 6 i_req_data[26]
port 89 nsew signal input
rlabel metal2 s 47712 99600 47768 100000 6 i_req_data[27]
port 90 nsew signal input
rlabel metal2 s 47936 99600 47992 100000 6 i_req_data[28]
port 91 nsew signal input
rlabel metal2 s 48160 99600 48216 100000 6 i_req_data[29]
port 92 nsew signal input
rlabel metal2 s 12096 99600 12152 100000 6 i_req_data[2]
port 93 nsew signal input
rlabel metal2 s 48384 99600 48440 100000 6 i_req_data[30]
port 94 nsew signal input
rlabel metal2 s 48608 99600 48664 100000 6 i_req_data[31]
port 95 nsew signal input
rlabel metal2 s 14784 99600 14840 100000 6 i_req_data[3]
port 96 nsew signal input
rlabel metal2 s 17472 99600 17528 100000 6 i_req_data[4]
port 97 nsew signal input
rlabel metal2 s 20160 99600 20216 100000 6 i_req_data[5]
port 98 nsew signal input
rlabel metal2 s 22848 99600 22904 100000 6 i_req_data[6]
port 99 nsew signal input
rlabel metal2 s 25536 99600 25592 100000 6 i_req_data[7]
port 100 nsew signal input
rlabel metal2 s 28224 99600 28280 100000 6 i_req_data[8]
port 101 nsew signal input
rlabel metal2 s 30464 99600 30520 100000 6 i_req_data[9]
port 102 nsew signal input
rlabel metal2 s 2688 99600 2744 100000 6 i_req_data_valid
port 103 nsew signal input
rlabel metal2 s 2912 99600 2968 100000 6 i_rst
port 104 nsew signal input
rlabel metal2 s 3136 99600 3192 100000 6 o_c_data_page
port 105 nsew signal output
rlabel metal2 s 3360 99600 3416 100000 6 o_c_instr_long
port 106 nsew signal output
rlabel metal2 s 3584 99600 3640 100000 6 o_c_instr_page
port 107 nsew signal output
rlabel metal2 s 3808 99600 3864 100000 6 o_icache_flush
port 108 nsew signal output
rlabel metal2 s 6496 99600 6552 100000 6 o_instr_long_addr[0]
port 109 nsew signal output
rlabel metal2 s 9408 99600 9464 100000 6 o_instr_long_addr[1]
port 110 nsew signal output
rlabel metal2 s 12320 99600 12376 100000 6 o_instr_long_addr[2]
port 111 nsew signal output
rlabel metal2 s 15008 99600 15064 100000 6 o_instr_long_addr[3]
port 112 nsew signal output
rlabel metal2 s 17696 99600 17752 100000 6 o_instr_long_addr[4]
port 113 nsew signal output
rlabel metal2 s 20384 99600 20440 100000 6 o_instr_long_addr[5]
port 114 nsew signal output
rlabel metal2 s 23072 99600 23128 100000 6 o_instr_long_addr[6]
port 115 nsew signal output
rlabel metal2 s 25760 99600 25816 100000 6 o_instr_long_addr[7]
port 116 nsew signal output
rlabel metal2 s 6720 99600 6776 100000 6 o_mem_addr[0]
port 117 nsew signal output
rlabel metal2 s 32928 99600 32984 100000 6 o_mem_addr[10]
port 118 nsew signal output
rlabel metal2 s 35168 99600 35224 100000 6 o_mem_addr[11]
port 119 nsew signal output
rlabel metal2 s 37408 99600 37464 100000 6 o_mem_addr[12]
port 120 nsew signal output
rlabel metal2 s 39648 99600 39704 100000 6 o_mem_addr[13]
port 121 nsew signal output
rlabel metal2 s 41888 99600 41944 100000 6 o_mem_addr[14]
port 122 nsew signal output
rlabel metal2 s 44128 99600 44184 100000 6 o_mem_addr[15]
port 123 nsew signal output
rlabel metal2 s 9632 99600 9688 100000 6 o_mem_addr[1]
port 124 nsew signal output
rlabel metal2 s 12544 99600 12600 100000 6 o_mem_addr[2]
port 125 nsew signal output
rlabel metal2 s 15232 99600 15288 100000 6 o_mem_addr[3]
port 126 nsew signal output
rlabel metal2 s 17920 99600 17976 100000 6 o_mem_addr[4]
port 127 nsew signal output
rlabel metal2 s 20608 99600 20664 100000 6 o_mem_addr[5]
port 128 nsew signal output
rlabel metal2 s 23296 99600 23352 100000 6 o_mem_addr[6]
port 129 nsew signal output
rlabel metal2 s 25984 99600 26040 100000 6 o_mem_addr[7]
port 130 nsew signal output
rlabel metal2 s 28448 99600 28504 100000 6 o_mem_addr[8]
port 131 nsew signal output
rlabel metal2 s 30688 99600 30744 100000 6 o_mem_addr[9]
port 132 nsew signal output
rlabel metal2 s 6944 99600 7000 100000 6 o_mem_addr_high[0]
port 133 nsew signal output
rlabel metal2 s 9856 99600 9912 100000 6 o_mem_addr_high[1]
port 134 nsew signal output
rlabel metal2 s 12768 99600 12824 100000 6 o_mem_addr_high[2]
port 135 nsew signal output
rlabel metal2 s 15456 99600 15512 100000 6 o_mem_addr_high[3]
port 136 nsew signal output
rlabel metal2 s 18144 99600 18200 100000 6 o_mem_addr_high[4]
port 137 nsew signal output
rlabel metal2 s 20832 99600 20888 100000 6 o_mem_addr_high[5]
port 138 nsew signal output
rlabel metal2 s 23520 99600 23576 100000 6 o_mem_addr_high[6]
port 139 nsew signal output
rlabel metal2 s 26208 99600 26264 100000 6 o_mem_addr_high[7]
port 140 nsew signal output
rlabel metal2 s 7168 99600 7224 100000 6 o_mem_data[0]
port 141 nsew signal output
rlabel metal2 s 33152 99600 33208 100000 6 o_mem_data[10]
port 142 nsew signal output
rlabel metal2 s 35392 99600 35448 100000 6 o_mem_data[11]
port 143 nsew signal output
rlabel metal2 s 37632 99600 37688 100000 6 o_mem_data[12]
port 144 nsew signal output
rlabel metal2 s 39872 99600 39928 100000 6 o_mem_data[13]
port 145 nsew signal output
rlabel metal2 s 42112 99600 42168 100000 6 o_mem_data[14]
port 146 nsew signal output
rlabel metal2 s 44352 99600 44408 100000 6 o_mem_data[15]
port 147 nsew signal output
rlabel metal2 s 10080 99600 10136 100000 6 o_mem_data[1]
port 148 nsew signal output
rlabel metal2 s 12992 99600 13048 100000 6 o_mem_data[2]
port 149 nsew signal output
rlabel metal2 s 15680 99600 15736 100000 6 o_mem_data[3]
port 150 nsew signal output
rlabel metal2 s 18368 99600 18424 100000 6 o_mem_data[4]
port 151 nsew signal output
rlabel metal2 s 21056 99600 21112 100000 6 o_mem_data[5]
port 152 nsew signal output
rlabel metal2 s 23744 99600 23800 100000 6 o_mem_data[6]
port 153 nsew signal output
rlabel metal2 s 26432 99600 26488 100000 6 o_mem_data[7]
port 154 nsew signal output
rlabel metal2 s 28672 99600 28728 100000 6 o_mem_data[8]
port 155 nsew signal output
rlabel metal2 s 30912 99600 30968 100000 6 o_mem_data[9]
port 156 nsew signal output
rlabel metal2 s 4032 99600 4088 100000 6 o_mem_long
port 157 nsew signal output
rlabel metal2 s 4256 99600 4312 100000 6 o_mem_req
port 158 nsew signal output
rlabel metal2 s 7392 99600 7448 100000 6 o_mem_sel[0]
port 159 nsew signal output
rlabel metal2 s 10304 99600 10360 100000 6 o_mem_sel[1]
port 160 nsew signal output
rlabel metal2 s 4480 99600 4536 100000 6 o_mem_we
port 161 nsew signal output
rlabel metal2 s 4704 99600 4760 100000 6 o_req_active
port 162 nsew signal output
rlabel metal2 s 7616 99600 7672 100000 6 o_req_addr[0]
port 163 nsew signal output
rlabel metal2 s 33376 99600 33432 100000 6 o_req_addr[10]
port 164 nsew signal output
rlabel metal2 s 35616 99600 35672 100000 6 o_req_addr[11]
port 165 nsew signal output
rlabel metal2 s 37856 99600 37912 100000 6 o_req_addr[12]
port 166 nsew signal output
rlabel metal2 s 40096 99600 40152 100000 6 o_req_addr[13]
port 167 nsew signal output
rlabel metal2 s 42336 99600 42392 100000 6 o_req_addr[14]
port 168 nsew signal output
rlabel metal2 s 44576 99600 44632 100000 6 o_req_addr[15]
port 169 nsew signal output
rlabel metal2 s 10528 99600 10584 100000 6 o_req_addr[1]
port 170 nsew signal output
rlabel metal2 s 13216 99600 13272 100000 6 o_req_addr[2]
port 171 nsew signal output
rlabel metal2 s 15904 99600 15960 100000 6 o_req_addr[3]
port 172 nsew signal output
rlabel metal2 s 18592 99600 18648 100000 6 o_req_addr[4]
port 173 nsew signal output
rlabel metal2 s 21280 99600 21336 100000 6 o_req_addr[5]
port 174 nsew signal output
rlabel metal2 s 23968 99600 24024 100000 6 o_req_addr[6]
port 175 nsew signal output
rlabel metal2 s 26656 99600 26712 100000 6 o_req_addr[7]
port 176 nsew signal output
rlabel metal2 s 28896 99600 28952 100000 6 o_req_addr[8]
port 177 nsew signal output
rlabel metal2 s 31136 99600 31192 100000 6 o_req_addr[9]
port 178 nsew signal output
rlabel metal2 s 4928 99600 4984 100000 6 o_req_ppl_submit
port 179 nsew signal output
rlabel metal2 s 7840 99600 7896 100000 6 sr_bus_addr[0]
port 180 nsew signal output
rlabel metal2 s 33600 99600 33656 100000 6 sr_bus_addr[10]
port 181 nsew signal output
rlabel metal2 s 35840 99600 35896 100000 6 sr_bus_addr[11]
port 182 nsew signal output
rlabel metal2 s 38080 99600 38136 100000 6 sr_bus_addr[12]
port 183 nsew signal output
rlabel metal2 s 40320 99600 40376 100000 6 sr_bus_addr[13]
port 184 nsew signal output
rlabel metal2 s 42560 99600 42616 100000 6 sr_bus_addr[14]
port 185 nsew signal output
rlabel metal2 s 44800 99600 44856 100000 6 sr_bus_addr[15]
port 186 nsew signal output
rlabel metal2 s 10752 99600 10808 100000 6 sr_bus_addr[1]
port 187 nsew signal output
rlabel metal2 s 13440 99600 13496 100000 6 sr_bus_addr[2]
port 188 nsew signal output
rlabel metal2 s 16128 99600 16184 100000 6 sr_bus_addr[3]
port 189 nsew signal output
rlabel metal2 s 18816 99600 18872 100000 6 sr_bus_addr[4]
port 190 nsew signal output
rlabel metal2 s 21504 99600 21560 100000 6 sr_bus_addr[5]
port 191 nsew signal output
rlabel metal2 s 24192 99600 24248 100000 6 sr_bus_addr[6]
port 192 nsew signal output
rlabel metal2 s 26880 99600 26936 100000 6 sr_bus_addr[7]
port 193 nsew signal output
rlabel metal2 s 29120 99600 29176 100000 6 sr_bus_addr[8]
port 194 nsew signal output
rlabel metal2 s 31360 99600 31416 100000 6 sr_bus_addr[9]
port 195 nsew signal output
rlabel metal2 s 8064 99600 8120 100000 6 sr_bus_data_o[0]
port 196 nsew signal output
rlabel metal2 s 33824 99600 33880 100000 6 sr_bus_data_o[10]
port 197 nsew signal output
rlabel metal2 s 36064 99600 36120 100000 6 sr_bus_data_o[11]
port 198 nsew signal output
rlabel metal2 s 38304 99600 38360 100000 6 sr_bus_data_o[12]
port 199 nsew signal output
rlabel metal2 s 40544 99600 40600 100000 6 sr_bus_data_o[13]
port 200 nsew signal output
rlabel metal2 s 42784 99600 42840 100000 6 sr_bus_data_o[14]
port 201 nsew signal output
rlabel metal2 s 45024 99600 45080 100000 6 sr_bus_data_o[15]
port 202 nsew signal output
rlabel metal2 s 10976 99600 11032 100000 6 sr_bus_data_o[1]
port 203 nsew signal output
rlabel metal2 s 13664 99600 13720 100000 6 sr_bus_data_o[2]
port 204 nsew signal output
rlabel metal2 s 16352 99600 16408 100000 6 sr_bus_data_o[3]
port 205 nsew signal output
rlabel metal2 s 19040 99600 19096 100000 6 sr_bus_data_o[4]
port 206 nsew signal output
rlabel metal2 s 21728 99600 21784 100000 6 sr_bus_data_o[5]
port 207 nsew signal output
rlabel metal2 s 24416 99600 24472 100000 6 sr_bus_data_o[6]
port 208 nsew signal output
rlabel metal2 s 27104 99600 27160 100000 6 sr_bus_data_o[7]
port 209 nsew signal output
rlabel metal2 s 29344 99600 29400 100000 6 sr_bus_data_o[8]
port 210 nsew signal output
rlabel metal2 s 31584 99600 31640 100000 6 sr_bus_data_o[9]
port 211 nsew signal output
rlabel metal2 s 5152 99600 5208 100000 6 sr_bus_we
port 212 nsew signal output
rlabel metal4 s 2224 1538 2384 98422 6 vccd1
port 213 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 98422 6 vccd1
port 213 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 98422 6 vccd1
port 213 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 98422 6 vccd1
port 213 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 98422 6 vssd1
port 214 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 98422 6 vssd1
port 214 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 98422 6 vssd1
port 214 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 50000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12912216
string GDS_FILE /home/piotro/caravel_user_project/openlane/core1/runs/23_11_12_10_40/results/signoff/core1.magic.gds
string GDS_START 592214
<< end >>

