// This is the unpowered netlist.
module interconnect_inner (c0_clk,
    c0_disable,
    c0_i_irq,
    c0_i_mc_core_int,
    c0_i_mem_ack,
    c0_i_mem_exception,
    c0_i_req_data_valid,
    c0_o_c_data_page,
    c0_o_c_instr_long,
    c0_o_c_instr_page,
    c0_o_icache_flush,
    c0_o_mem_long_mode,
    c0_o_mem_req,
    c0_o_mem_we,
    c0_o_req_active,
    c0_o_req_ppl_submit,
    c0_rst,
    c0_sr_bus_we,
    c1_clk,
    c1_disable,
    c1_i_irq,
    c1_i_mc_core_int,
    c1_i_mem_ack,
    c1_i_mem_exception,
    c1_i_req_data_valid,
    c1_o_c_data_page,
    c1_o_c_instr_long,
    c1_o_c_instr_page,
    c1_o_icache_flush,
    c1_o_mem_long_mode,
    c1_o_mem_req,
    c1_o_mem_we,
    c1_o_req_active,
    c1_o_req_ppl_submit,
    c1_rst,
    c1_sr_bus_we,
    core_clock,
    core_reset,
    dcache_clk,
    dcache_mem_ack,
    dcache_mem_cache_enable,
    dcache_mem_exception,
    dcache_mem_req,
    dcache_mem_we,
    dcache_rst,
    dcache_wb_4_burst,
    dcache_wb_ack,
    dcache_wb_cyc,
    dcache_wb_err,
    dcache_wb_stb,
    dcache_wb_we,
    ic0_clk,
    ic0_mem_ack,
    ic0_mem_cache_flush,
    ic0_mem_ppl_submit,
    ic0_mem_req,
    ic0_rst,
    ic0_wb_ack,
    ic0_wb_cyc,
    ic0_wb_err,
    ic0_wb_stb,
    ic0_wb_we,
    ic1_clk,
    ic1_mem_ack,
    ic1_mem_cache_flush,
    ic1_mem_ppl_submit,
    ic1_mem_req,
    ic1_rst,
    ic1_wb_ack,
    ic1_wb_cyc,
    ic1_wb_err,
    ic1_wb_stb,
    ic1_wb_we,
    inner_disable,
    inner_embed_mode,
    inner_ext_irq,
    inner_wb_4_burst,
    inner_wb_8_burst,
    inner_wb_ack,
    inner_wb_cyc,
    inner_wb_err,
    inner_wb_stb,
    inner_wb_we,
    c0_dbg_pc,
    c0_dbg_r0,
    c0_i_core_int_sreg,
    c0_i_mem_data,
    c0_i_req_data,
    c0_o_instr_long_addr,
    c0_o_mem_addr,
    c0_o_mem_data,
    c0_o_mem_high_addr,
    c0_o_mem_sel,
    c0_o_req_addr,
    c0_sr_bus_addr,
    c0_sr_bus_data_o,
    c1_dbg_pc,
    c1_dbg_r0,
    c1_i_core_int_sreg,
    c1_i_mem_data,
    c1_i_req_data,
    c1_o_instr_long_addr,
    c1_o_mem_addr,
    c1_o_mem_data,
    c1_o_mem_high_addr,
    c1_o_mem_sel,
    c1_o_req_addr,
    c1_sr_bus_addr,
    c1_sr_bus_data_o,
    dcache_mem_addr,
    dcache_mem_i_data,
    dcache_mem_o_data,
    dcache_mem_sel,
    dcache_wb_adr,
    dcache_wb_i_dat,
    dcache_wb_o_dat,
    dcache_wb_sel,
    ic0_mem_addr,
    ic0_mem_data,
    ic0_wb_adr,
    ic0_wb_i_dat,
    ic0_wb_sel,
    ic1_mem_addr,
    ic1_mem_data,
    ic1_wb_adr,
    ic1_wb_i_dat,
    ic1_wb_sel,
    inner_wb_adr,
    inner_wb_i_dat,
    inner_wb_o_dat,
    inner_wb_sel);
 output c0_clk;
 output c0_disable;
 output c0_i_irq;
 output c0_i_mc_core_int;
 output c0_i_mem_ack;
 output c0_i_mem_exception;
 output c0_i_req_data_valid;
 input c0_o_c_data_page;
 input c0_o_c_instr_long;
 input c0_o_c_instr_page;
 input c0_o_icache_flush;
 input c0_o_mem_long_mode;
 input c0_o_mem_req;
 input c0_o_mem_we;
 input c0_o_req_active;
 input c0_o_req_ppl_submit;
 output c0_rst;
 input c0_sr_bus_we;
 output c1_clk;
 output c1_disable;
 output c1_i_irq;
 output c1_i_mc_core_int;
 output c1_i_mem_ack;
 output c1_i_mem_exception;
 output c1_i_req_data_valid;
 input c1_o_c_data_page;
 input c1_o_c_instr_long;
 input c1_o_c_instr_page;
 input c1_o_icache_flush;
 input c1_o_mem_long_mode;
 input c1_o_mem_req;
 input c1_o_mem_we;
 input c1_o_req_active;
 input c1_o_req_ppl_submit;
 output c1_rst;
 input c1_sr_bus_we;
 input core_clock;
 input core_reset;
 output dcache_clk;
 input dcache_mem_ack;
 output dcache_mem_cache_enable;
 input dcache_mem_exception;
 output dcache_mem_req;
 output dcache_mem_we;
 output dcache_rst;
 input dcache_wb_4_burst;
 output dcache_wb_ack;
 input dcache_wb_cyc;
 output dcache_wb_err;
 input dcache_wb_stb;
 input dcache_wb_we;
 output ic0_clk;
 input ic0_mem_ack;
 output ic0_mem_cache_flush;
 output ic0_mem_ppl_submit;
 output ic0_mem_req;
 output ic0_rst;
 output ic0_wb_ack;
 input ic0_wb_cyc;
 output ic0_wb_err;
 input ic0_wb_stb;
 input ic0_wb_we;
 output ic1_clk;
 input ic1_mem_ack;
 output ic1_mem_cache_flush;
 output ic1_mem_ppl_submit;
 output ic1_mem_req;
 output ic1_rst;
 output ic1_wb_ack;
 input ic1_wb_cyc;
 output ic1_wb_err;
 input ic1_wb_stb;
 input ic1_wb_we;
 input inner_disable;
 input inner_embed_mode;
 input inner_ext_irq;
 output inner_wb_4_burst;
 output inner_wb_8_burst;
 input inner_wb_ack;
 output inner_wb_cyc;
 input inner_wb_err;
 output inner_wb_stb;
 output inner_wb_we;
 input [15:0] c0_dbg_pc;
 input [15:0] c0_dbg_r0;
 output [15:0] c0_i_core_int_sreg;
 output [15:0] c0_i_mem_data;
 output [31:0] c0_i_req_data;
 input [7:0] c0_o_instr_long_addr;
 input [15:0] c0_o_mem_addr;
 input [15:0] c0_o_mem_data;
 input [7:0] c0_o_mem_high_addr;
 input [1:0] c0_o_mem_sel;
 input [15:0] c0_o_req_addr;
 input [15:0] c0_sr_bus_addr;
 input [15:0] c0_sr_bus_data_o;
 input [15:0] c1_dbg_pc;
 input [15:0] c1_dbg_r0;
 output [15:0] c1_i_core_int_sreg;
 output [15:0] c1_i_mem_data;
 output [31:0] c1_i_req_data;
 input [7:0] c1_o_instr_long_addr;
 input [15:0] c1_o_mem_addr;
 input [15:0] c1_o_mem_data;
 input [7:0] c1_o_mem_high_addr;
 input [1:0] c1_o_mem_sel;
 input [15:0] c1_o_req_addr;
 input [15:0] c1_sr_bus_addr;
 input [15:0] c1_sr_bus_data_o;
 output [23:0] dcache_mem_addr;
 output [15:0] dcache_mem_i_data;
 input [15:0] dcache_mem_o_data;
 output [1:0] dcache_mem_sel;
 input [23:0] dcache_wb_adr;
 output [15:0] dcache_wb_i_dat;
 input [15:0] dcache_wb_o_dat;
 input [1:0] dcache_wb_sel;
 output [15:0] ic0_mem_addr;
 input [31:0] ic0_mem_data;
 input [15:0] ic0_wb_adr;
 output [15:0] ic0_wb_i_dat;
 input [1:0] ic0_wb_sel;
 output [15:0] ic1_mem_addr;
 input [31:0] ic1_mem_data;
 input [15:0] ic1_wb_adr;
 output [15:0] ic1_wb_i_dat;
 input [1:0] ic1_wb_sel;
 output [23:0] inner_wb_adr;
 input [15:0] inner_wb_i_dat;
 output [15:0] inner_wb_o_dat;
 output [1:0] inner_wb_sel;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire clknet_leaf_0_core_clock;
 wire \dmmu0.long_off_reg[0] ;
 wire \dmmu0.long_off_reg[1] ;
 wire \dmmu0.long_off_reg[2] ;
 wire \dmmu0.long_off_reg[3] ;
 wire \dmmu0.long_off_reg[4] ;
 wire \dmmu0.long_off_reg[5] ;
 wire \dmmu0.long_off_reg[6] ;
 wire \dmmu0.long_off_reg[7] ;
 wire \dmmu0.page_table[0][0] ;
 wire \dmmu0.page_table[0][10] ;
 wire \dmmu0.page_table[0][11] ;
 wire \dmmu0.page_table[0][12] ;
 wire \dmmu0.page_table[0][1] ;
 wire \dmmu0.page_table[0][2] ;
 wire \dmmu0.page_table[0][3] ;
 wire \dmmu0.page_table[0][4] ;
 wire \dmmu0.page_table[0][5] ;
 wire \dmmu0.page_table[0][6] ;
 wire \dmmu0.page_table[0][7] ;
 wire \dmmu0.page_table[0][8] ;
 wire \dmmu0.page_table[0][9] ;
 wire \dmmu0.page_table[10][0] ;
 wire \dmmu0.page_table[10][10] ;
 wire \dmmu0.page_table[10][11] ;
 wire \dmmu0.page_table[10][12] ;
 wire \dmmu0.page_table[10][1] ;
 wire \dmmu0.page_table[10][2] ;
 wire \dmmu0.page_table[10][3] ;
 wire \dmmu0.page_table[10][4] ;
 wire \dmmu0.page_table[10][5] ;
 wire \dmmu0.page_table[10][6] ;
 wire \dmmu0.page_table[10][7] ;
 wire \dmmu0.page_table[10][8] ;
 wire \dmmu0.page_table[10][9] ;
 wire \dmmu0.page_table[11][0] ;
 wire \dmmu0.page_table[11][10] ;
 wire \dmmu0.page_table[11][11] ;
 wire \dmmu0.page_table[11][12] ;
 wire \dmmu0.page_table[11][1] ;
 wire \dmmu0.page_table[11][2] ;
 wire \dmmu0.page_table[11][3] ;
 wire \dmmu0.page_table[11][4] ;
 wire \dmmu0.page_table[11][5] ;
 wire \dmmu0.page_table[11][6] ;
 wire \dmmu0.page_table[11][7] ;
 wire \dmmu0.page_table[11][8] ;
 wire \dmmu0.page_table[11][9] ;
 wire \dmmu0.page_table[12][0] ;
 wire \dmmu0.page_table[12][10] ;
 wire \dmmu0.page_table[12][11] ;
 wire \dmmu0.page_table[12][12] ;
 wire \dmmu0.page_table[12][1] ;
 wire \dmmu0.page_table[12][2] ;
 wire \dmmu0.page_table[12][3] ;
 wire \dmmu0.page_table[12][4] ;
 wire \dmmu0.page_table[12][5] ;
 wire \dmmu0.page_table[12][6] ;
 wire \dmmu0.page_table[12][7] ;
 wire \dmmu0.page_table[12][8] ;
 wire \dmmu0.page_table[12][9] ;
 wire \dmmu0.page_table[13][0] ;
 wire \dmmu0.page_table[13][10] ;
 wire \dmmu0.page_table[13][11] ;
 wire \dmmu0.page_table[13][12] ;
 wire \dmmu0.page_table[13][1] ;
 wire \dmmu0.page_table[13][2] ;
 wire \dmmu0.page_table[13][3] ;
 wire \dmmu0.page_table[13][4] ;
 wire \dmmu0.page_table[13][5] ;
 wire \dmmu0.page_table[13][6] ;
 wire \dmmu0.page_table[13][7] ;
 wire \dmmu0.page_table[13][8] ;
 wire \dmmu0.page_table[13][9] ;
 wire \dmmu0.page_table[14][0] ;
 wire \dmmu0.page_table[14][10] ;
 wire \dmmu0.page_table[14][11] ;
 wire \dmmu0.page_table[14][12] ;
 wire \dmmu0.page_table[14][1] ;
 wire \dmmu0.page_table[14][2] ;
 wire \dmmu0.page_table[14][3] ;
 wire \dmmu0.page_table[14][4] ;
 wire \dmmu0.page_table[14][5] ;
 wire \dmmu0.page_table[14][6] ;
 wire \dmmu0.page_table[14][7] ;
 wire \dmmu0.page_table[14][8] ;
 wire \dmmu0.page_table[14][9] ;
 wire \dmmu0.page_table[15][0] ;
 wire \dmmu0.page_table[15][10] ;
 wire \dmmu0.page_table[15][11] ;
 wire \dmmu0.page_table[15][12] ;
 wire \dmmu0.page_table[15][1] ;
 wire \dmmu0.page_table[15][2] ;
 wire \dmmu0.page_table[15][3] ;
 wire \dmmu0.page_table[15][4] ;
 wire \dmmu0.page_table[15][5] ;
 wire \dmmu0.page_table[15][6] ;
 wire \dmmu0.page_table[15][7] ;
 wire \dmmu0.page_table[15][8] ;
 wire \dmmu0.page_table[15][9] ;
 wire \dmmu0.page_table[1][0] ;
 wire \dmmu0.page_table[1][10] ;
 wire \dmmu0.page_table[1][11] ;
 wire \dmmu0.page_table[1][12] ;
 wire \dmmu0.page_table[1][1] ;
 wire \dmmu0.page_table[1][2] ;
 wire \dmmu0.page_table[1][3] ;
 wire \dmmu0.page_table[1][4] ;
 wire \dmmu0.page_table[1][5] ;
 wire \dmmu0.page_table[1][6] ;
 wire \dmmu0.page_table[1][7] ;
 wire \dmmu0.page_table[1][8] ;
 wire \dmmu0.page_table[1][9] ;
 wire \dmmu0.page_table[2][0] ;
 wire \dmmu0.page_table[2][10] ;
 wire \dmmu0.page_table[2][11] ;
 wire \dmmu0.page_table[2][12] ;
 wire \dmmu0.page_table[2][1] ;
 wire \dmmu0.page_table[2][2] ;
 wire \dmmu0.page_table[2][3] ;
 wire \dmmu0.page_table[2][4] ;
 wire \dmmu0.page_table[2][5] ;
 wire \dmmu0.page_table[2][6] ;
 wire \dmmu0.page_table[2][7] ;
 wire \dmmu0.page_table[2][8] ;
 wire \dmmu0.page_table[2][9] ;
 wire \dmmu0.page_table[3][0] ;
 wire \dmmu0.page_table[3][10] ;
 wire \dmmu0.page_table[3][11] ;
 wire \dmmu0.page_table[3][12] ;
 wire \dmmu0.page_table[3][1] ;
 wire \dmmu0.page_table[3][2] ;
 wire \dmmu0.page_table[3][3] ;
 wire \dmmu0.page_table[3][4] ;
 wire \dmmu0.page_table[3][5] ;
 wire \dmmu0.page_table[3][6] ;
 wire \dmmu0.page_table[3][7] ;
 wire \dmmu0.page_table[3][8] ;
 wire \dmmu0.page_table[3][9] ;
 wire \dmmu0.page_table[4][0] ;
 wire \dmmu0.page_table[4][10] ;
 wire \dmmu0.page_table[4][11] ;
 wire \dmmu0.page_table[4][12] ;
 wire \dmmu0.page_table[4][1] ;
 wire \dmmu0.page_table[4][2] ;
 wire \dmmu0.page_table[4][3] ;
 wire \dmmu0.page_table[4][4] ;
 wire \dmmu0.page_table[4][5] ;
 wire \dmmu0.page_table[4][6] ;
 wire \dmmu0.page_table[4][7] ;
 wire \dmmu0.page_table[4][8] ;
 wire \dmmu0.page_table[4][9] ;
 wire \dmmu0.page_table[5][0] ;
 wire \dmmu0.page_table[5][10] ;
 wire \dmmu0.page_table[5][11] ;
 wire \dmmu0.page_table[5][12] ;
 wire \dmmu0.page_table[5][1] ;
 wire \dmmu0.page_table[5][2] ;
 wire \dmmu0.page_table[5][3] ;
 wire \dmmu0.page_table[5][4] ;
 wire \dmmu0.page_table[5][5] ;
 wire \dmmu0.page_table[5][6] ;
 wire \dmmu0.page_table[5][7] ;
 wire \dmmu0.page_table[5][8] ;
 wire \dmmu0.page_table[5][9] ;
 wire \dmmu0.page_table[6][0] ;
 wire \dmmu0.page_table[6][10] ;
 wire \dmmu0.page_table[6][11] ;
 wire \dmmu0.page_table[6][12] ;
 wire \dmmu0.page_table[6][1] ;
 wire \dmmu0.page_table[6][2] ;
 wire \dmmu0.page_table[6][3] ;
 wire \dmmu0.page_table[6][4] ;
 wire \dmmu0.page_table[6][5] ;
 wire \dmmu0.page_table[6][6] ;
 wire \dmmu0.page_table[6][7] ;
 wire \dmmu0.page_table[6][8] ;
 wire \dmmu0.page_table[6][9] ;
 wire \dmmu0.page_table[7][0] ;
 wire \dmmu0.page_table[7][10] ;
 wire \dmmu0.page_table[7][11] ;
 wire \dmmu0.page_table[7][12] ;
 wire \dmmu0.page_table[7][1] ;
 wire \dmmu0.page_table[7][2] ;
 wire \dmmu0.page_table[7][3] ;
 wire \dmmu0.page_table[7][4] ;
 wire \dmmu0.page_table[7][5] ;
 wire \dmmu0.page_table[7][6] ;
 wire \dmmu0.page_table[7][7] ;
 wire \dmmu0.page_table[7][8] ;
 wire \dmmu0.page_table[7][9] ;
 wire \dmmu0.page_table[8][0] ;
 wire \dmmu0.page_table[8][10] ;
 wire \dmmu0.page_table[8][11] ;
 wire \dmmu0.page_table[8][12] ;
 wire \dmmu0.page_table[8][1] ;
 wire \dmmu0.page_table[8][2] ;
 wire \dmmu0.page_table[8][3] ;
 wire \dmmu0.page_table[8][4] ;
 wire \dmmu0.page_table[8][5] ;
 wire \dmmu0.page_table[8][6] ;
 wire \dmmu0.page_table[8][7] ;
 wire \dmmu0.page_table[8][8] ;
 wire \dmmu0.page_table[8][9] ;
 wire \dmmu0.page_table[9][0] ;
 wire \dmmu0.page_table[9][10] ;
 wire \dmmu0.page_table[9][11] ;
 wire \dmmu0.page_table[9][12] ;
 wire \dmmu0.page_table[9][1] ;
 wire \dmmu0.page_table[9][2] ;
 wire \dmmu0.page_table[9][3] ;
 wire \dmmu0.page_table[9][4] ;
 wire \dmmu0.page_table[9][5] ;
 wire \dmmu0.page_table[9][6] ;
 wire \dmmu0.page_table[9][7] ;
 wire \dmmu0.page_table[9][8] ;
 wire \dmmu0.page_table[9][9] ;
 wire \dmmu1.long_off_reg[0] ;
 wire \dmmu1.long_off_reg[1] ;
 wire \dmmu1.long_off_reg[2] ;
 wire \dmmu1.long_off_reg[3] ;
 wire \dmmu1.long_off_reg[4] ;
 wire \dmmu1.long_off_reg[5] ;
 wire \dmmu1.long_off_reg[6] ;
 wire \dmmu1.long_off_reg[7] ;
 wire \dmmu1.page_table[0][0] ;
 wire \dmmu1.page_table[0][10] ;
 wire \dmmu1.page_table[0][11] ;
 wire \dmmu1.page_table[0][12] ;
 wire \dmmu1.page_table[0][1] ;
 wire \dmmu1.page_table[0][2] ;
 wire \dmmu1.page_table[0][3] ;
 wire \dmmu1.page_table[0][4] ;
 wire \dmmu1.page_table[0][5] ;
 wire \dmmu1.page_table[0][6] ;
 wire \dmmu1.page_table[0][7] ;
 wire \dmmu1.page_table[0][8] ;
 wire \dmmu1.page_table[0][9] ;
 wire \dmmu1.page_table[10][0] ;
 wire \dmmu1.page_table[10][10] ;
 wire \dmmu1.page_table[10][11] ;
 wire \dmmu1.page_table[10][12] ;
 wire \dmmu1.page_table[10][1] ;
 wire \dmmu1.page_table[10][2] ;
 wire \dmmu1.page_table[10][3] ;
 wire \dmmu1.page_table[10][4] ;
 wire \dmmu1.page_table[10][5] ;
 wire \dmmu1.page_table[10][6] ;
 wire \dmmu1.page_table[10][7] ;
 wire \dmmu1.page_table[10][8] ;
 wire \dmmu1.page_table[10][9] ;
 wire \dmmu1.page_table[11][0] ;
 wire \dmmu1.page_table[11][10] ;
 wire \dmmu1.page_table[11][11] ;
 wire \dmmu1.page_table[11][12] ;
 wire \dmmu1.page_table[11][1] ;
 wire \dmmu1.page_table[11][2] ;
 wire \dmmu1.page_table[11][3] ;
 wire \dmmu1.page_table[11][4] ;
 wire \dmmu1.page_table[11][5] ;
 wire \dmmu1.page_table[11][6] ;
 wire \dmmu1.page_table[11][7] ;
 wire \dmmu1.page_table[11][8] ;
 wire \dmmu1.page_table[11][9] ;
 wire \dmmu1.page_table[12][0] ;
 wire \dmmu1.page_table[12][10] ;
 wire \dmmu1.page_table[12][11] ;
 wire \dmmu1.page_table[12][12] ;
 wire \dmmu1.page_table[12][1] ;
 wire \dmmu1.page_table[12][2] ;
 wire \dmmu1.page_table[12][3] ;
 wire \dmmu1.page_table[12][4] ;
 wire \dmmu1.page_table[12][5] ;
 wire \dmmu1.page_table[12][6] ;
 wire \dmmu1.page_table[12][7] ;
 wire \dmmu1.page_table[12][8] ;
 wire \dmmu1.page_table[12][9] ;
 wire \dmmu1.page_table[13][0] ;
 wire \dmmu1.page_table[13][10] ;
 wire \dmmu1.page_table[13][11] ;
 wire \dmmu1.page_table[13][12] ;
 wire \dmmu1.page_table[13][1] ;
 wire \dmmu1.page_table[13][2] ;
 wire \dmmu1.page_table[13][3] ;
 wire \dmmu1.page_table[13][4] ;
 wire \dmmu1.page_table[13][5] ;
 wire \dmmu1.page_table[13][6] ;
 wire \dmmu1.page_table[13][7] ;
 wire \dmmu1.page_table[13][8] ;
 wire \dmmu1.page_table[13][9] ;
 wire \dmmu1.page_table[14][0] ;
 wire \dmmu1.page_table[14][10] ;
 wire \dmmu1.page_table[14][11] ;
 wire \dmmu1.page_table[14][12] ;
 wire \dmmu1.page_table[14][1] ;
 wire \dmmu1.page_table[14][2] ;
 wire \dmmu1.page_table[14][3] ;
 wire \dmmu1.page_table[14][4] ;
 wire \dmmu1.page_table[14][5] ;
 wire \dmmu1.page_table[14][6] ;
 wire \dmmu1.page_table[14][7] ;
 wire \dmmu1.page_table[14][8] ;
 wire \dmmu1.page_table[14][9] ;
 wire \dmmu1.page_table[15][0] ;
 wire \dmmu1.page_table[15][10] ;
 wire \dmmu1.page_table[15][11] ;
 wire \dmmu1.page_table[15][12] ;
 wire \dmmu1.page_table[15][1] ;
 wire \dmmu1.page_table[15][2] ;
 wire \dmmu1.page_table[15][3] ;
 wire \dmmu1.page_table[15][4] ;
 wire \dmmu1.page_table[15][5] ;
 wire \dmmu1.page_table[15][6] ;
 wire \dmmu1.page_table[15][7] ;
 wire \dmmu1.page_table[15][8] ;
 wire \dmmu1.page_table[15][9] ;
 wire \dmmu1.page_table[1][0] ;
 wire \dmmu1.page_table[1][10] ;
 wire \dmmu1.page_table[1][11] ;
 wire \dmmu1.page_table[1][12] ;
 wire \dmmu1.page_table[1][1] ;
 wire \dmmu1.page_table[1][2] ;
 wire \dmmu1.page_table[1][3] ;
 wire \dmmu1.page_table[1][4] ;
 wire \dmmu1.page_table[1][5] ;
 wire \dmmu1.page_table[1][6] ;
 wire \dmmu1.page_table[1][7] ;
 wire \dmmu1.page_table[1][8] ;
 wire \dmmu1.page_table[1][9] ;
 wire \dmmu1.page_table[2][0] ;
 wire \dmmu1.page_table[2][10] ;
 wire \dmmu1.page_table[2][11] ;
 wire \dmmu1.page_table[2][12] ;
 wire \dmmu1.page_table[2][1] ;
 wire \dmmu1.page_table[2][2] ;
 wire \dmmu1.page_table[2][3] ;
 wire \dmmu1.page_table[2][4] ;
 wire \dmmu1.page_table[2][5] ;
 wire \dmmu1.page_table[2][6] ;
 wire \dmmu1.page_table[2][7] ;
 wire \dmmu1.page_table[2][8] ;
 wire \dmmu1.page_table[2][9] ;
 wire \dmmu1.page_table[3][0] ;
 wire \dmmu1.page_table[3][10] ;
 wire \dmmu1.page_table[3][11] ;
 wire \dmmu1.page_table[3][12] ;
 wire \dmmu1.page_table[3][1] ;
 wire \dmmu1.page_table[3][2] ;
 wire \dmmu1.page_table[3][3] ;
 wire \dmmu1.page_table[3][4] ;
 wire \dmmu1.page_table[3][5] ;
 wire \dmmu1.page_table[3][6] ;
 wire \dmmu1.page_table[3][7] ;
 wire \dmmu1.page_table[3][8] ;
 wire \dmmu1.page_table[3][9] ;
 wire \dmmu1.page_table[4][0] ;
 wire \dmmu1.page_table[4][10] ;
 wire \dmmu1.page_table[4][11] ;
 wire \dmmu1.page_table[4][12] ;
 wire \dmmu1.page_table[4][1] ;
 wire \dmmu1.page_table[4][2] ;
 wire \dmmu1.page_table[4][3] ;
 wire \dmmu1.page_table[4][4] ;
 wire \dmmu1.page_table[4][5] ;
 wire \dmmu1.page_table[4][6] ;
 wire \dmmu1.page_table[4][7] ;
 wire \dmmu1.page_table[4][8] ;
 wire \dmmu1.page_table[4][9] ;
 wire \dmmu1.page_table[5][0] ;
 wire \dmmu1.page_table[5][10] ;
 wire \dmmu1.page_table[5][11] ;
 wire \dmmu1.page_table[5][12] ;
 wire \dmmu1.page_table[5][1] ;
 wire \dmmu1.page_table[5][2] ;
 wire \dmmu1.page_table[5][3] ;
 wire \dmmu1.page_table[5][4] ;
 wire \dmmu1.page_table[5][5] ;
 wire \dmmu1.page_table[5][6] ;
 wire \dmmu1.page_table[5][7] ;
 wire \dmmu1.page_table[5][8] ;
 wire \dmmu1.page_table[5][9] ;
 wire \dmmu1.page_table[6][0] ;
 wire \dmmu1.page_table[6][10] ;
 wire \dmmu1.page_table[6][11] ;
 wire \dmmu1.page_table[6][12] ;
 wire \dmmu1.page_table[6][1] ;
 wire \dmmu1.page_table[6][2] ;
 wire \dmmu1.page_table[6][3] ;
 wire \dmmu1.page_table[6][4] ;
 wire \dmmu1.page_table[6][5] ;
 wire \dmmu1.page_table[6][6] ;
 wire \dmmu1.page_table[6][7] ;
 wire \dmmu1.page_table[6][8] ;
 wire \dmmu1.page_table[6][9] ;
 wire \dmmu1.page_table[7][0] ;
 wire \dmmu1.page_table[7][10] ;
 wire \dmmu1.page_table[7][11] ;
 wire \dmmu1.page_table[7][12] ;
 wire \dmmu1.page_table[7][1] ;
 wire \dmmu1.page_table[7][2] ;
 wire \dmmu1.page_table[7][3] ;
 wire \dmmu1.page_table[7][4] ;
 wire \dmmu1.page_table[7][5] ;
 wire \dmmu1.page_table[7][6] ;
 wire \dmmu1.page_table[7][7] ;
 wire \dmmu1.page_table[7][8] ;
 wire \dmmu1.page_table[7][9] ;
 wire \dmmu1.page_table[8][0] ;
 wire \dmmu1.page_table[8][10] ;
 wire \dmmu1.page_table[8][11] ;
 wire \dmmu1.page_table[8][12] ;
 wire \dmmu1.page_table[8][1] ;
 wire \dmmu1.page_table[8][2] ;
 wire \dmmu1.page_table[8][3] ;
 wire \dmmu1.page_table[8][4] ;
 wire \dmmu1.page_table[8][5] ;
 wire \dmmu1.page_table[8][6] ;
 wire \dmmu1.page_table[8][7] ;
 wire \dmmu1.page_table[8][8] ;
 wire \dmmu1.page_table[8][9] ;
 wire \dmmu1.page_table[9][0] ;
 wire \dmmu1.page_table[9][10] ;
 wire \dmmu1.page_table[9][11] ;
 wire \dmmu1.page_table[9][12] ;
 wire \dmmu1.page_table[9][1] ;
 wire \dmmu1.page_table[9][2] ;
 wire \dmmu1.page_table[9][3] ;
 wire \dmmu1.page_table[9][4] ;
 wire \dmmu1.page_table[9][5] ;
 wire \dmmu1.page_table[9][6] ;
 wire \dmmu1.page_table[9][7] ;
 wire \dmmu1.page_table[9][8] ;
 wire \dmmu1.page_table[9][9] ;
 wire \icache_arbiter.o_sel_sig ;
 wire \icore_sregs.c1_disable ;
 wire \immu_0.high_addr_off[0] ;
 wire \immu_0.high_addr_off[1] ;
 wire \immu_0.high_addr_off[2] ;
 wire \immu_0.high_addr_off[3] ;
 wire \immu_0.high_addr_off[4] ;
 wire \immu_0.high_addr_off[5] ;
 wire \immu_0.high_addr_off[6] ;
 wire \immu_0.high_addr_off[7] ;
 wire \immu_0.page_table[0][0] ;
 wire \immu_0.page_table[0][10] ;
 wire \immu_0.page_table[0][1] ;
 wire \immu_0.page_table[0][2] ;
 wire \immu_0.page_table[0][3] ;
 wire \immu_0.page_table[0][4] ;
 wire \immu_0.page_table[0][5] ;
 wire \immu_0.page_table[0][6] ;
 wire \immu_0.page_table[0][7] ;
 wire \immu_0.page_table[0][8] ;
 wire \immu_0.page_table[0][9] ;
 wire \immu_0.page_table[10][0] ;
 wire \immu_0.page_table[10][10] ;
 wire \immu_0.page_table[10][1] ;
 wire \immu_0.page_table[10][2] ;
 wire \immu_0.page_table[10][3] ;
 wire \immu_0.page_table[10][4] ;
 wire \immu_0.page_table[10][5] ;
 wire \immu_0.page_table[10][6] ;
 wire \immu_0.page_table[10][7] ;
 wire \immu_0.page_table[10][8] ;
 wire \immu_0.page_table[10][9] ;
 wire \immu_0.page_table[11][0] ;
 wire \immu_0.page_table[11][10] ;
 wire \immu_0.page_table[11][1] ;
 wire \immu_0.page_table[11][2] ;
 wire \immu_0.page_table[11][3] ;
 wire \immu_0.page_table[11][4] ;
 wire \immu_0.page_table[11][5] ;
 wire \immu_0.page_table[11][6] ;
 wire \immu_0.page_table[11][7] ;
 wire \immu_0.page_table[11][8] ;
 wire \immu_0.page_table[11][9] ;
 wire \immu_0.page_table[12][0] ;
 wire \immu_0.page_table[12][10] ;
 wire \immu_0.page_table[12][1] ;
 wire \immu_0.page_table[12][2] ;
 wire \immu_0.page_table[12][3] ;
 wire \immu_0.page_table[12][4] ;
 wire \immu_0.page_table[12][5] ;
 wire \immu_0.page_table[12][6] ;
 wire \immu_0.page_table[12][7] ;
 wire \immu_0.page_table[12][8] ;
 wire \immu_0.page_table[12][9] ;
 wire \immu_0.page_table[13][0] ;
 wire \immu_0.page_table[13][10] ;
 wire \immu_0.page_table[13][1] ;
 wire \immu_0.page_table[13][2] ;
 wire \immu_0.page_table[13][3] ;
 wire \immu_0.page_table[13][4] ;
 wire \immu_0.page_table[13][5] ;
 wire \immu_0.page_table[13][6] ;
 wire \immu_0.page_table[13][7] ;
 wire \immu_0.page_table[13][8] ;
 wire \immu_0.page_table[13][9] ;
 wire \immu_0.page_table[14][0] ;
 wire \immu_0.page_table[14][10] ;
 wire \immu_0.page_table[14][1] ;
 wire \immu_0.page_table[14][2] ;
 wire \immu_0.page_table[14][3] ;
 wire \immu_0.page_table[14][4] ;
 wire \immu_0.page_table[14][5] ;
 wire \immu_0.page_table[14][6] ;
 wire \immu_0.page_table[14][7] ;
 wire \immu_0.page_table[14][8] ;
 wire \immu_0.page_table[14][9] ;
 wire \immu_0.page_table[15][0] ;
 wire \immu_0.page_table[15][10] ;
 wire \immu_0.page_table[15][1] ;
 wire \immu_0.page_table[15][2] ;
 wire \immu_0.page_table[15][3] ;
 wire \immu_0.page_table[15][4] ;
 wire \immu_0.page_table[15][5] ;
 wire \immu_0.page_table[15][6] ;
 wire \immu_0.page_table[15][7] ;
 wire \immu_0.page_table[15][8] ;
 wire \immu_0.page_table[15][9] ;
 wire \immu_0.page_table[1][0] ;
 wire \immu_0.page_table[1][10] ;
 wire \immu_0.page_table[1][1] ;
 wire \immu_0.page_table[1][2] ;
 wire \immu_0.page_table[1][3] ;
 wire \immu_0.page_table[1][4] ;
 wire \immu_0.page_table[1][5] ;
 wire \immu_0.page_table[1][6] ;
 wire \immu_0.page_table[1][7] ;
 wire \immu_0.page_table[1][8] ;
 wire \immu_0.page_table[1][9] ;
 wire \immu_0.page_table[2][0] ;
 wire \immu_0.page_table[2][10] ;
 wire \immu_0.page_table[2][1] ;
 wire \immu_0.page_table[2][2] ;
 wire \immu_0.page_table[2][3] ;
 wire \immu_0.page_table[2][4] ;
 wire \immu_0.page_table[2][5] ;
 wire \immu_0.page_table[2][6] ;
 wire \immu_0.page_table[2][7] ;
 wire \immu_0.page_table[2][8] ;
 wire \immu_0.page_table[2][9] ;
 wire \immu_0.page_table[3][0] ;
 wire \immu_0.page_table[3][10] ;
 wire \immu_0.page_table[3][1] ;
 wire \immu_0.page_table[3][2] ;
 wire \immu_0.page_table[3][3] ;
 wire \immu_0.page_table[3][4] ;
 wire \immu_0.page_table[3][5] ;
 wire \immu_0.page_table[3][6] ;
 wire \immu_0.page_table[3][7] ;
 wire \immu_0.page_table[3][8] ;
 wire \immu_0.page_table[3][9] ;
 wire \immu_0.page_table[4][0] ;
 wire \immu_0.page_table[4][10] ;
 wire \immu_0.page_table[4][1] ;
 wire \immu_0.page_table[4][2] ;
 wire \immu_0.page_table[4][3] ;
 wire \immu_0.page_table[4][4] ;
 wire \immu_0.page_table[4][5] ;
 wire \immu_0.page_table[4][6] ;
 wire \immu_0.page_table[4][7] ;
 wire \immu_0.page_table[4][8] ;
 wire \immu_0.page_table[4][9] ;
 wire \immu_0.page_table[5][0] ;
 wire \immu_0.page_table[5][10] ;
 wire \immu_0.page_table[5][1] ;
 wire \immu_0.page_table[5][2] ;
 wire \immu_0.page_table[5][3] ;
 wire \immu_0.page_table[5][4] ;
 wire \immu_0.page_table[5][5] ;
 wire \immu_0.page_table[5][6] ;
 wire \immu_0.page_table[5][7] ;
 wire \immu_0.page_table[5][8] ;
 wire \immu_0.page_table[5][9] ;
 wire \immu_0.page_table[6][0] ;
 wire \immu_0.page_table[6][10] ;
 wire \immu_0.page_table[6][1] ;
 wire \immu_0.page_table[6][2] ;
 wire \immu_0.page_table[6][3] ;
 wire \immu_0.page_table[6][4] ;
 wire \immu_0.page_table[6][5] ;
 wire \immu_0.page_table[6][6] ;
 wire \immu_0.page_table[6][7] ;
 wire \immu_0.page_table[6][8] ;
 wire \immu_0.page_table[6][9] ;
 wire \immu_0.page_table[7][0] ;
 wire \immu_0.page_table[7][10] ;
 wire \immu_0.page_table[7][1] ;
 wire \immu_0.page_table[7][2] ;
 wire \immu_0.page_table[7][3] ;
 wire \immu_0.page_table[7][4] ;
 wire \immu_0.page_table[7][5] ;
 wire \immu_0.page_table[7][6] ;
 wire \immu_0.page_table[7][7] ;
 wire \immu_0.page_table[7][8] ;
 wire \immu_0.page_table[7][9] ;
 wire \immu_0.page_table[8][0] ;
 wire \immu_0.page_table[8][10] ;
 wire \immu_0.page_table[8][1] ;
 wire \immu_0.page_table[8][2] ;
 wire \immu_0.page_table[8][3] ;
 wire \immu_0.page_table[8][4] ;
 wire \immu_0.page_table[8][5] ;
 wire \immu_0.page_table[8][6] ;
 wire \immu_0.page_table[8][7] ;
 wire \immu_0.page_table[8][8] ;
 wire \immu_0.page_table[8][9] ;
 wire \immu_0.page_table[9][0] ;
 wire \immu_0.page_table[9][10] ;
 wire \immu_0.page_table[9][1] ;
 wire \immu_0.page_table[9][2] ;
 wire \immu_0.page_table[9][3] ;
 wire \immu_0.page_table[9][4] ;
 wire \immu_0.page_table[9][5] ;
 wire \immu_0.page_table[9][6] ;
 wire \immu_0.page_table[9][7] ;
 wire \immu_0.page_table[9][8] ;
 wire \immu_0.page_table[9][9] ;
 wire \immu_1.high_addr_off[0] ;
 wire \immu_1.high_addr_off[1] ;
 wire \immu_1.high_addr_off[2] ;
 wire \immu_1.high_addr_off[3] ;
 wire \immu_1.high_addr_off[4] ;
 wire \immu_1.high_addr_off[5] ;
 wire \immu_1.high_addr_off[6] ;
 wire \immu_1.high_addr_off[7] ;
 wire \immu_1.page_table[0][0] ;
 wire \immu_1.page_table[0][10] ;
 wire \immu_1.page_table[0][1] ;
 wire \immu_1.page_table[0][2] ;
 wire \immu_1.page_table[0][3] ;
 wire \immu_1.page_table[0][4] ;
 wire \immu_1.page_table[0][5] ;
 wire \immu_1.page_table[0][6] ;
 wire \immu_1.page_table[0][7] ;
 wire \immu_1.page_table[0][8] ;
 wire \immu_1.page_table[0][9] ;
 wire \immu_1.page_table[10][0] ;
 wire \immu_1.page_table[10][10] ;
 wire \immu_1.page_table[10][1] ;
 wire \immu_1.page_table[10][2] ;
 wire \immu_1.page_table[10][3] ;
 wire \immu_1.page_table[10][4] ;
 wire \immu_1.page_table[10][5] ;
 wire \immu_1.page_table[10][6] ;
 wire \immu_1.page_table[10][7] ;
 wire \immu_1.page_table[10][8] ;
 wire \immu_1.page_table[10][9] ;
 wire \immu_1.page_table[11][0] ;
 wire \immu_1.page_table[11][10] ;
 wire \immu_1.page_table[11][1] ;
 wire \immu_1.page_table[11][2] ;
 wire \immu_1.page_table[11][3] ;
 wire \immu_1.page_table[11][4] ;
 wire \immu_1.page_table[11][5] ;
 wire \immu_1.page_table[11][6] ;
 wire \immu_1.page_table[11][7] ;
 wire \immu_1.page_table[11][8] ;
 wire \immu_1.page_table[11][9] ;
 wire \immu_1.page_table[12][0] ;
 wire \immu_1.page_table[12][10] ;
 wire \immu_1.page_table[12][1] ;
 wire \immu_1.page_table[12][2] ;
 wire \immu_1.page_table[12][3] ;
 wire \immu_1.page_table[12][4] ;
 wire \immu_1.page_table[12][5] ;
 wire \immu_1.page_table[12][6] ;
 wire \immu_1.page_table[12][7] ;
 wire \immu_1.page_table[12][8] ;
 wire \immu_1.page_table[12][9] ;
 wire \immu_1.page_table[13][0] ;
 wire \immu_1.page_table[13][10] ;
 wire \immu_1.page_table[13][1] ;
 wire \immu_1.page_table[13][2] ;
 wire \immu_1.page_table[13][3] ;
 wire \immu_1.page_table[13][4] ;
 wire \immu_1.page_table[13][5] ;
 wire \immu_1.page_table[13][6] ;
 wire \immu_1.page_table[13][7] ;
 wire \immu_1.page_table[13][8] ;
 wire \immu_1.page_table[13][9] ;
 wire \immu_1.page_table[14][0] ;
 wire \immu_1.page_table[14][10] ;
 wire \immu_1.page_table[14][1] ;
 wire \immu_1.page_table[14][2] ;
 wire \immu_1.page_table[14][3] ;
 wire \immu_1.page_table[14][4] ;
 wire \immu_1.page_table[14][5] ;
 wire \immu_1.page_table[14][6] ;
 wire \immu_1.page_table[14][7] ;
 wire \immu_1.page_table[14][8] ;
 wire \immu_1.page_table[14][9] ;
 wire \immu_1.page_table[15][0] ;
 wire \immu_1.page_table[15][10] ;
 wire \immu_1.page_table[15][1] ;
 wire \immu_1.page_table[15][2] ;
 wire \immu_1.page_table[15][3] ;
 wire \immu_1.page_table[15][4] ;
 wire \immu_1.page_table[15][5] ;
 wire \immu_1.page_table[15][6] ;
 wire \immu_1.page_table[15][7] ;
 wire \immu_1.page_table[15][8] ;
 wire \immu_1.page_table[15][9] ;
 wire \immu_1.page_table[1][0] ;
 wire \immu_1.page_table[1][10] ;
 wire \immu_1.page_table[1][1] ;
 wire \immu_1.page_table[1][2] ;
 wire \immu_1.page_table[1][3] ;
 wire \immu_1.page_table[1][4] ;
 wire \immu_1.page_table[1][5] ;
 wire \immu_1.page_table[1][6] ;
 wire \immu_1.page_table[1][7] ;
 wire \immu_1.page_table[1][8] ;
 wire \immu_1.page_table[1][9] ;
 wire \immu_1.page_table[2][0] ;
 wire \immu_1.page_table[2][10] ;
 wire \immu_1.page_table[2][1] ;
 wire \immu_1.page_table[2][2] ;
 wire \immu_1.page_table[2][3] ;
 wire \immu_1.page_table[2][4] ;
 wire \immu_1.page_table[2][5] ;
 wire \immu_1.page_table[2][6] ;
 wire \immu_1.page_table[2][7] ;
 wire \immu_1.page_table[2][8] ;
 wire \immu_1.page_table[2][9] ;
 wire \immu_1.page_table[3][0] ;
 wire \immu_1.page_table[3][10] ;
 wire \immu_1.page_table[3][1] ;
 wire \immu_1.page_table[3][2] ;
 wire \immu_1.page_table[3][3] ;
 wire \immu_1.page_table[3][4] ;
 wire \immu_1.page_table[3][5] ;
 wire \immu_1.page_table[3][6] ;
 wire \immu_1.page_table[3][7] ;
 wire \immu_1.page_table[3][8] ;
 wire \immu_1.page_table[3][9] ;
 wire \immu_1.page_table[4][0] ;
 wire \immu_1.page_table[4][10] ;
 wire \immu_1.page_table[4][1] ;
 wire \immu_1.page_table[4][2] ;
 wire \immu_1.page_table[4][3] ;
 wire \immu_1.page_table[4][4] ;
 wire \immu_1.page_table[4][5] ;
 wire \immu_1.page_table[4][6] ;
 wire \immu_1.page_table[4][7] ;
 wire \immu_1.page_table[4][8] ;
 wire \immu_1.page_table[4][9] ;
 wire \immu_1.page_table[5][0] ;
 wire \immu_1.page_table[5][10] ;
 wire \immu_1.page_table[5][1] ;
 wire \immu_1.page_table[5][2] ;
 wire \immu_1.page_table[5][3] ;
 wire \immu_1.page_table[5][4] ;
 wire \immu_1.page_table[5][5] ;
 wire \immu_1.page_table[5][6] ;
 wire \immu_1.page_table[5][7] ;
 wire \immu_1.page_table[5][8] ;
 wire \immu_1.page_table[5][9] ;
 wire \immu_1.page_table[6][0] ;
 wire \immu_1.page_table[6][10] ;
 wire \immu_1.page_table[6][1] ;
 wire \immu_1.page_table[6][2] ;
 wire \immu_1.page_table[6][3] ;
 wire \immu_1.page_table[6][4] ;
 wire \immu_1.page_table[6][5] ;
 wire \immu_1.page_table[6][6] ;
 wire \immu_1.page_table[6][7] ;
 wire \immu_1.page_table[6][8] ;
 wire \immu_1.page_table[6][9] ;
 wire \immu_1.page_table[7][0] ;
 wire \immu_1.page_table[7][10] ;
 wire \immu_1.page_table[7][1] ;
 wire \immu_1.page_table[7][2] ;
 wire \immu_1.page_table[7][3] ;
 wire \immu_1.page_table[7][4] ;
 wire \immu_1.page_table[7][5] ;
 wire \immu_1.page_table[7][6] ;
 wire \immu_1.page_table[7][7] ;
 wire \immu_1.page_table[7][8] ;
 wire \immu_1.page_table[7][9] ;
 wire \immu_1.page_table[8][0] ;
 wire \immu_1.page_table[8][10] ;
 wire \immu_1.page_table[8][1] ;
 wire \immu_1.page_table[8][2] ;
 wire \immu_1.page_table[8][3] ;
 wire \immu_1.page_table[8][4] ;
 wire \immu_1.page_table[8][5] ;
 wire \immu_1.page_table[8][6] ;
 wire \immu_1.page_table[8][7] ;
 wire \immu_1.page_table[8][8] ;
 wire \immu_1.page_table[8][9] ;
 wire \immu_1.page_table[9][0] ;
 wire \immu_1.page_table[9][10] ;
 wire \immu_1.page_table[9][1] ;
 wire \immu_1.page_table[9][2] ;
 wire \immu_1.page_table[9][3] ;
 wire \immu_1.page_table[9][4] ;
 wire \immu_1.page_table[9][5] ;
 wire \immu_1.page_table[9][6] ;
 wire \immu_1.page_table[9][7] ;
 wire \immu_1.page_table[9][8] ;
 wire \immu_1.page_table[9][9] ;
 wire \inner_wb_arbiter.o_sel_sig ;
 wire \mem_dcache_arb.req0_pending ;
 wire \mem_dcache_arb.req1_pending ;
 wire \mem_dcache_arb.select ;
 wire \mem_dcache_arb.transfer_active ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire clknet_leaf_1_core_clock;
 wire clknet_leaf_2_core_clock;
 wire clknet_leaf_3_core_clock;
 wire clknet_leaf_4_core_clock;
 wire clknet_leaf_5_core_clock;
 wire clknet_leaf_6_core_clock;
 wire clknet_leaf_7_core_clock;
 wire clknet_leaf_8_core_clock;
 wire clknet_leaf_9_core_clock;
 wire clknet_leaf_10_core_clock;
 wire clknet_leaf_11_core_clock;
 wire clknet_leaf_12_core_clock;
 wire clknet_leaf_13_core_clock;
 wire clknet_leaf_14_core_clock;
 wire clknet_leaf_15_core_clock;
 wire clknet_leaf_16_core_clock;
 wire clknet_leaf_17_core_clock;
 wire clknet_leaf_18_core_clock;
 wire clknet_leaf_19_core_clock;
 wire clknet_leaf_20_core_clock;
 wire clknet_leaf_21_core_clock;
 wire clknet_leaf_22_core_clock;
 wire clknet_leaf_23_core_clock;
 wire clknet_leaf_24_core_clock;
 wire clknet_leaf_25_core_clock;
 wire clknet_leaf_26_core_clock;
 wire clknet_leaf_27_core_clock;
 wire clknet_leaf_28_core_clock;
 wire clknet_leaf_29_core_clock;
 wire clknet_leaf_30_core_clock;
 wire clknet_leaf_31_core_clock;
 wire clknet_leaf_32_core_clock;
 wire clknet_leaf_33_core_clock;
 wire clknet_leaf_34_core_clock;
 wire clknet_leaf_35_core_clock;
 wire clknet_leaf_36_core_clock;
 wire clknet_leaf_37_core_clock;
 wire clknet_leaf_38_core_clock;
 wire clknet_leaf_39_core_clock;
 wire clknet_leaf_40_core_clock;
 wire clknet_leaf_41_core_clock;
 wire clknet_leaf_42_core_clock;
 wire clknet_leaf_43_core_clock;
 wire clknet_leaf_44_core_clock;
 wire clknet_leaf_45_core_clock;
 wire clknet_leaf_46_core_clock;
 wire clknet_leaf_47_core_clock;
 wire clknet_leaf_48_core_clock;
 wire clknet_leaf_49_core_clock;
 wire clknet_leaf_50_core_clock;
 wire clknet_leaf_51_core_clock;
 wire clknet_leaf_53_core_clock;
 wire clknet_leaf_54_core_clock;
 wire clknet_leaf_55_core_clock;
 wire clknet_leaf_56_core_clock;
 wire clknet_leaf_57_core_clock;
 wire clknet_leaf_58_core_clock;
 wire clknet_leaf_59_core_clock;
 wire clknet_leaf_60_core_clock;
 wire clknet_leaf_61_core_clock;
 wire clknet_leaf_62_core_clock;
 wire clknet_leaf_63_core_clock;
 wire clknet_leaf_66_core_clock;
 wire clknet_leaf_67_core_clock;
 wire clknet_leaf_68_core_clock;
 wire clknet_leaf_69_core_clock;
 wire clknet_leaf_70_core_clock;
 wire clknet_leaf_71_core_clock;
 wire clknet_leaf_72_core_clock;
 wire clknet_leaf_73_core_clock;
 wire clknet_leaf_74_core_clock;
 wire clknet_leaf_75_core_clock;
 wire clknet_leaf_76_core_clock;
 wire clknet_leaf_77_core_clock;
 wire clknet_leaf_78_core_clock;
 wire clknet_leaf_79_core_clock;
 wire clknet_leaf_80_core_clock;
 wire clknet_leaf_81_core_clock;
 wire clknet_leaf_82_core_clock;
 wire clknet_leaf_83_core_clock;
 wire clknet_leaf_84_core_clock;
 wire clknet_leaf_85_core_clock;
 wire clknet_leaf_86_core_clock;
 wire clknet_leaf_87_core_clock;
 wire clknet_leaf_88_core_clock;
 wire clknet_leaf_89_core_clock;
 wire clknet_leaf_90_core_clock;
 wire clknet_leaf_91_core_clock;
 wire clknet_leaf_92_core_clock;
 wire clknet_leaf_93_core_clock;
 wire clknet_0_core_clock;
 wire clknet_1_0_0_core_clock;
 wire clknet_1_0_1_core_clock;
 wire clknet_1_1_0_core_clock;
 wire clknet_1_1_1_core_clock;
 wire clknet_2_0_0_core_clock;
 wire clknet_2_1_0_core_clock;
 wire clknet_2_2_0_core_clock;
 wire clknet_2_3_0_core_clock;
 wire clknet_3_0_0_core_clock;
 wire clknet_3_1_0_core_clock;
 wire clknet_3_2_0_core_clock;
 wire clknet_3_3_0_core_clock;
 wire clknet_3_4_0_core_clock;
 wire clknet_3_5_0_core_clock;
 wire clknet_3_6_0_core_clock;
 wire clknet_3_7_0_core_clock;
 wire clknet_opt_1_0_core_clock;
 wire clknet_opt_2_0_core_clock;
 wire clknet_opt_2_1_core_clock;

 sky130_fd_sc_hd__nor2_2 _3184_ (.A(\mem_dcache_arb.req0_pending ),
    .B(net54),
    .Y(_0809_));
 sky130_fd_sc_hd__nor2_4 _3185_ (.A(\mem_dcache_arb.req1_pending ),
    .B(net159),
    .Y(_0810_));
 sky130_fd_sc_hd__a21oi_4 _3186_ (.A1(_0809_),
    .A2(_0810_),
    .B1(\mem_dcache_arb.transfer_active ),
    .Y(net562));
 sky130_fd_sc_hd__inv_6 _3187_ (.A(\inner_wb_arbiter.o_sel_sig ),
    .Y(_0811_));
 sky130_fd_sc_hd__buf_12 _3188_ (.A(_0811_),
    .X(net664));
 sky130_fd_sc_hd__buf_6 _3189_ (.A(\icache_arbiter.o_sel_sig ),
    .X(_0812_));
 sky130_fd_sc_hd__inv_6 _3190_ (.A(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__and3_1 _3191_ (.A(net664),
    .B(_0813_),
    .C(net387),
    .X(_0814_));
 sky130_fd_sc_hd__clkbuf_1 _3192_ (.A(_0814_),
    .X(net606));
 sky130_fd_sc_hd__and3_1 _3193_ (.A(net664),
    .B(_0813_),
    .C(net388),
    .X(_0815_));
 sky130_fd_sc_hd__clkbuf_1 _3194_ (.A(_0815_),
    .X(net607));
 sky130_fd_sc_hd__nor2_1 _3195_ (.A(\mem_dcache_arb.select ),
    .B(_0810_),
    .Y(_0816_));
 sky130_fd_sc_hd__or3_2 _3196_ (.A(\mem_dcache_arb.transfer_active ),
    .B(_0809_),
    .C(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__o21a_2 _3197_ (.A1(\mem_dcache_arb.select ),
    .A2(net562),
    .B1(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__clkbuf_4 _3198_ (.A(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__and2_1 _3199_ (.A(net214),
    .B(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__clkbuf_1 _3200_ (.A(_0820_),
    .X(net469));
 sky130_fd_sc_hd__and2_1 _3201_ (.A(net221),
    .B(_0819_),
    .X(_0821_));
 sky130_fd_sc_hd__clkbuf_1 _3202_ (.A(_0821_),
    .X(net476));
 sky130_fd_sc_hd__and2_1 _3203_ (.A(net222),
    .B(_0819_),
    .X(_0822_));
 sky130_fd_sc_hd__clkbuf_1 _3204_ (.A(_0822_),
    .X(net477));
 sky130_fd_sc_hd__and2_1 _3205_ (.A(net223),
    .B(_0819_),
    .X(_0823_));
 sky130_fd_sc_hd__clkbuf_1 _3206_ (.A(_0823_),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_2 _3207_ (.A(_0818_),
    .X(_0824_));
 sky130_fd_sc_hd__and2_1 _3208_ (.A(net224),
    .B(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__clkbuf_1 _3209_ (.A(_0825_),
    .X(net479));
 sky130_fd_sc_hd__and2_1 _3210_ (.A(net225),
    .B(_0824_),
    .X(_0826_));
 sky130_fd_sc_hd__clkbuf_1 _3211_ (.A(_0826_),
    .X(net480));
 sky130_fd_sc_hd__and2_1 _3212_ (.A(net226),
    .B(_0824_),
    .X(_0827_));
 sky130_fd_sc_hd__clkbuf_1 _3213_ (.A(_0827_),
    .X(net481));
 sky130_fd_sc_hd__and2_1 _3214_ (.A(net227),
    .B(_0824_),
    .X(_0828_));
 sky130_fd_sc_hd__clkbuf_1 _3215_ (.A(_0828_),
    .X(net482));
 sky130_fd_sc_hd__and2_1 _3216_ (.A(net228),
    .B(_0824_),
    .X(_0829_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3217_ (.A(_0829_),
    .X(net483));
 sky130_fd_sc_hd__and2_1 _3218_ (.A(net229),
    .B(_0824_),
    .X(_0830_));
 sky130_fd_sc_hd__clkbuf_1 _3219_ (.A(_0830_),
    .X(net484));
 sky130_fd_sc_hd__and2_1 _3220_ (.A(net215),
    .B(_0824_),
    .X(_0831_));
 sky130_fd_sc_hd__clkbuf_1 _3221_ (.A(_0831_),
    .X(net470));
 sky130_fd_sc_hd__and2_1 _3222_ (.A(net216),
    .B(_0824_),
    .X(_0832_));
 sky130_fd_sc_hd__clkbuf_1 _3223_ (.A(_0832_),
    .X(net471));
 sky130_fd_sc_hd__and2_1 _3224_ (.A(net217),
    .B(_0824_),
    .X(_0833_));
 sky130_fd_sc_hd__clkbuf_1 _3225_ (.A(_0833_),
    .X(net472));
 sky130_fd_sc_hd__and2_1 _3226_ (.A(net218),
    .B(_0824_),
    .X(_0834_));
 sky130_fd_sc_hd__clkbuf_1 _3227_ (.A(_0834_),
    .X(net473));
 sky130_fd_sc_hd__buf_4 _3228_ (.A(_0818_),
    .X(_0835_));
 sky130_fd_sc_hd__and2_2 _3229_ (.A(net219),
    .B(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__clkbuf_1 _3230_ (.A(_0836_),
    .X(net474));
 sky130_fd_sc_hd__and2_2 _3231_ (.A(net220),
    .B(_0835_),
    .X(_0837_));
 sky130_fd_sc_hd__clkbuf_1 _3232_ (.A(_0837_),
    .X(net475));
 sky130_fd_sc_hd__o21ai_2 _3233_ (.A1(\mem_dcache_arb.select ),
    .A2(net562),
    .B1(_0817_),
    .Y(_0838_));
 sky130_fd_sc_hd__clkbuf_8 _3234_ (.A(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__buf_6 _3235_ (.A(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _3236_ (.A0(net162),
    .A1(net57),
    .S(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__clkbuf_1 _3237_ (.A(_0841_),
    .X(net565));
 sky130_fd_sc_hd__mux2_1 _3238_ (.A0(net118),
    .A1(net13),
    .S(_0840_),
    .X(_0842_));
 sky130_fd_sc_hd__clkbuf_1 _3239_ (.A(_0842_),
    .X(net521));
 sky130_fd_sc_hd__mux2_1 _3240_ (.A0(net125),
    .A1(net20),
    .S(_0840_),
    .X(_0843_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3241_ (.A(_0843_),
    .X(net532));
 sky130_fd_sc_hd__mux2_1 _3242_ (.A0(net126),
    .A1(net21),
    .S(_0840_),
    .X(_0844_));
 sky130_fd_sc_hd__clkbuf_1 _3243_ (.A(_0844_),
    .X(net537));
 sky130_fd_sc_hd__mux2_1 _3244_ (.A0(net127),
    .A1(net22),
    .S(_0840_),
    .X(_0845_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3245_ (.A(_0845_),
    .X(net538));
 sky130_fd_sc_hd__mux2_2 _3246_ (.A0(net128),
    .A1(net23),
    .S(_0840_),
    .X(_0846_));
 sky130_fd_sc_hd__clkbuf_1 _3247_ (.A(_0846_),
    .X(net539));
 sky130_fd_sc_hd__buf_4 _3248_ (.A(_0839_),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_2 _3249_ (.A0(net129),
    .A1(net24),
    .S(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__clkbuf_1 _3250_ (.A(_0848_),
    .X(net540));
 sky130_fd_sc_hd__mux2_2 _3251_ (.A0(net130),
    .A1(net25),
    .S(_0847_),
    .X(_0849_));
 sky130_fd_sc_hd__clkbuf_1 _3252_ (.A(_0849_),
    .X(net541));
 sky130_fd_sc_hd__mux2_2 _3253_ (.A0(net131),
    .A1(net26),
    .S(_0847_),
    .X(_0850_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3254_ (.A(_0850_),
    .X(net542));
 sky130_fd_sc_hd__mux2_2 _3255_ (.A0(net132),
    .A1(net27),
    .S(_0847_),
    .X(_0851_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3256_ (.A(_0851_),
    .X(net543));
 sky130_fd_sc_hd__mux2_2 _3257_ (.A0(net133),
    .A1(net28),
    .S(_0847_),
    .X(_0852_));
 sky130_fd_sc_hd__clkbuf_2 _3258_ (.A(_0852_),
    .X(net544));
 sky130_fd_sc_hd__mux2_2 _3259_ (.A0(net119),
    .A1(net14),
    .S(_0847_),
    .X(_0853_));
 sky130_fd_sc_hd__clkbuf_2 _3260_ (.A(_0853_),
    .X(net522));
 sky130_fd_sc_hd__buf_4 _3261_ (.A(net122),
    .X(_0854_));
 sky130_fd_sc_hd__buf_4 _3262_ (.A(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__buf_4 _3263_ (.A(net120),
    .X(_0856_));
 sky130_fd_sc_hd__buf_6 _3264_ (.A(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__buf_6 _3265_ (.A(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__clkbuf_4 _3266_ (.A(net121),
    .X(_0859_));
 sky130_fd_sc_hd__buf_4 _3267_ (.A(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__buf_4 _3268_ (.A(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__mux4_1 _3269_ (.A0(\dmmu1.page_table[12][0] ),
    .A1(\dmmu1.page_table[13][0] ),
    .A2(\dmmu1.page_table[14][0] ),
    .A3(\dmmu1.page_table[15][0] ),
    .S0(_0858_),
    .S1(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__clkbuf_4 _3270_ (.A(_0860_),
    .X(_0863_));
 sky130_fd_sc_hd__clkbuf_4 _3271_ (.A(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__buf_6 _3272_ (.A(_0857_),
    .X(_0865_));
 sky130_fd_sc_hd__mux2_1 _3273_ (.A0(\dmmu1.page_table[8][0] ),
    .A1(\dmmu1.page_table[9][0] ),
    .S(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__or2_1 _3274_ (.A(_0864_),
    .B(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__inv_2 _3275_ (.A(net121),
    .Y(_0868_));
 sky130_fd_sc_hd__clkbuf_8 _3276_ (.A(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__mux2_1 _3277_ (.A0(\dmmu1.page_table[10][0] ),
    .A1(\dmmu1.page_table[11][0] ),
    .S(_0858_),
    .X(_0870_));
 sky130_fd_sc_hd__inv_2 _3278_ (.A(net122),
    .Y(_0871_));
 sky130_fd_sc_hd__buf_4 _3279_ (.A(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__o21a_1 _3280_ (.A1(_0869_),
    .A2(_0870_),
    .B1(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__inv_6 _3281_ (.A(net123),
    .Y(_0874_));
 sky130_fd_sc_hd__a221o_1 _3282_ (.A1(_0855_),
    .A2(_0862_),
    .B1(_0867_),
    .B2(_0873_),
    .C1(_0874_),
    .X(_0875_));
 sky130_fd_sc_hd__or4_1 _3283_ (.A(net155),
    .B(net154),
    .C(net157),
    .D(net156),
    .X(_0876_));
 sky130_fd_sc_hd__or4_1 _3284_ (.A(net151),
    .B(net150),
    .C(net153),
    .D(net152),
    .X(_0877_));
 sky130_fd_sc_hd__or3_2 _3285_ (.A(net124),
    .B(_0876_),
    .C(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__nand2_4 _3286_ (.A(net158),
    .B(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__o21a_2 _3287_ (.A1(net106),
    .A2(net158),
    .B1(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__buf_4 _3288_ (.A(_0872_),
    .X(_0881_));
 sky130_fd_sc_hd__mux2_1 _3289_ (.A0(\dmmu1.page_table[0][0] ),
    .A1(\dmmu1.page_table[1][0] ),
    .S(_0865_),
    .X(_0882_));
 sky130_fd_sc_hd__or2_1 _3290_ (.A(_0864_),
    .B(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _3291_ (.A0(\dmmu1.page_table[2][0] ),
    .A1(\dmmu1.page_table[3][0] ),
    .S(_0865_),
    .X(_0884_));
 sky130_fd_sc_hd__or2_1 _3292_ (.A(_0869_),
    .B(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__mux4_1 _3293_ (.A0(\dmmu1.page_table[4][0] ),
    .A1(\dmmu1.page_table[5][0] ),
    .A2(\dmmu1.page_table[6][0] ),
    .A3(\dmmu1.page_table[7][0] ),
    .S0(_0865_),
    .S1(_0863_),
    .X(_0886_));
 sky130_fd_sc_hd__buf_4 _3294_ (.A(net123),
    .X(_0887_));
 sky130_fd_sc_hd__a21o_1 _3295_ (.A1(_0855_),
    .A2(_0886_),
    .B1(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__a31o_1 _3296_ (.A1(_0881_),
    .A2(_0883_),
    .A3(_0885_),
    .B1(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__and3_2 _3297_ (.A(_0875_),
    .B(_0880_),
    .C(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__buf_6 _3298_ (.A(_0857_),
    .X(_0891_));
 sky130_fd_sc_hd__buf_6 _3299_ (.A(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__o21ai_2 _3300_ (.A1(net106),
    .A2(net158),
    .B1(_0879_),
    .Y(_0893_));
 sky130_fd_sc_hd__a21o_1 _3301_ (.A1(_0892_),
    .A2(_0893_),
    .B1(_0840_),
    .X(_0894_));
 sky130_fd_sc_hd__buf_4 _3302_ (.A(net15),
    .X(_0895_));
 sky130_fd_sc_hd__buf_6 _3303_ (.A(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__buf_6 _3304_ (.A(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__buf_6 _3305_ (.A(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__buf_2 _3306_ (.A(net18),
    .X(_0899_));
 sky130_fd_sc_hd__buf_6 _3307_ (.A(_0896_),
    .X(_0900_));
 sky130_fd_sc_hd__clkbuf_4 _3308_ (.A(net16),
    .X(_0901_));
 sky130_fd_sc_hd__buf_4 _3309_ (.A(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__mux4_1 _3310_ (.A0(\dmmu0.page_table[0][0] ),
    .A1(\dmmu0.page_table[1][0] ),
    .A2(\dmmu0.page_table[2][0] ),
    .A3(\dmmu0.page_table[3][0] ),
    .S0(_0900_),
    .S1(_0902_),
    .X(_0903_));
 sky130_fd_sc_hd__mux4_1 _3311_ (.A0(\dmmu0.page_table[4][0] ),
    .A1(\dmmu0.page_table[5][0] ),
    .A2(\dmmu0.page_table[6][0] ),
    .A3(\dmmu0.page_table[7][0] ),
    .S0(_0900_),
    .S1(_0902_),
    .X(_0904_));
 sky130_fd_sc_hd__buf_4 _3312_ (.A(net17),
    .X(_0905_));
 sky130_fd_sc_hd__buf_4 _3313_ (.A(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_1 _3314_ (.A0(_0903_),
    .A1(_0904_),
    .S(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__inv_2 _3315_ (.A(net16),
    .Y(_0908_));
 sky130_fd_sc_hd__buf_4 _3316_ (.A(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__buf_6 _3317_ (.A(_0900_),
    .X(_0910_));
 sky130_fd_sc_hd__mux2_1 _3318_ (.A0(\dmmu0.page_table[14][0] ),
    .A1(\dmmu0.page_table[15][0] ),
    .S(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__clkbuf_8 _3319_ (.A(_0901_),
    .X(_0912_));
 sky130_fd_sc_hd__buf_4 _3320_ (.A(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _3321_ (.A0(\dmmu0.page_table[12][0] ),
    .A1(\dmmu0.page_table[13][0] ),
    .S(_0900_),
    .X(_0914_));
 sky130_fd_sc_hd__or2_1 _3322_ (.A(_0913_),
    .B(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__o211a_1 _3323_ (.A1(_0909_),
    .A2(_0911_),
    .B1(_0915_),
    .C1(_0906_),
    .X(_0916_));
 sky130_fd_sc_hd__clkinv_4 _3324_ (.A(net17),
    .Y(_0917_));
 sky130_fd_sc_hd__buf_4 _3325_ (.A(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__mux4_1 _3326_ (.A0(\dmmu0.page_table[8][0] ),
    .A1(\dmmu0.page_table[9][0] ),
    .A2(\dmmu0.page_table[10][0] ),
    .A3(\dmmu0.page_table[11][0] ),
    .S0(_0897_),
    .S1(_0902_),
    .X(_0919_));
 sky130_fd_sc_hd__inv_2 _3327_ (.A(net18),
    .Y(_0920_));
 sky130_fd_sc_hd__buf_4 _3328_ (.A(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__a21o_1 _3329_ (.A1(_0918_),
    .A2(_0919_),
    .B1(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__o22a_1 _3330_ (.A1(_0899_),
    .A2(_0907_),
    .B1(_0916_),
    .B2(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__or4_1 _3331_ (.A(net50),
    .B(net49),
    .C(net52),
    .D(net51),
    .X(_0924_));
 sky130_fd_sc_hd__or4_1 _3332_ (.A(net46),
    .B(net45),
    .C(net48),
    .D(net47),
    .X(_0925_));
 sky130_fd_sc_hd__or3_1 _3333_ (.A(net19),
    .B(_0924_),
    .C(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__and2_1 _3334_ (.A(net53),
    .B(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__nor2_2 _3335_ (.A(net1),
    .B(net53),
    .Y(_0928_));
 sky130_fd_sc_hd__nor2_4 _3336_ (.A(_0927_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__mux2_1 _3337_ (.A0(_0898_),
    .A1(_0923_),
    .S(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__o22a_2 _3338_ (.A1(_0890_),
    .A2(_0894_),
    .B1(_0930_),
    .B2(_0819_),
    .X(net523));
 sky130_fd_sc_hd__mux2_1 _3339_ (.A0(\dmmu1.page_table[14][1] ),
    .A1(\dmmu1.page_table[15][1] ),
    .S(_0865_),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_1 _3340_ (.A0(\dmmu1.page_table[12][1] ),
    .A1(\dmmu1.page_table[13][1] ),
    .S(_0857_),
    .X(_0932_));
 sky130_fd_sc_hd__or2_1 _3341_ (.A(_0863_),
    .B(_0932_),
    .X(_0933_));
 sky130_fd_sc_hd__o211a_1 _3342_ (.A1(_0869_),
    .A2(_0931_),
    .B1(_0933_),
    .C1(_0854_),
    .X(_0934_));
 sky130_fd_sc_hd__mux4_1 _3343_ (.A0(\dmmu1.page_table[8][1] ),
    .A1(\dmmu1.page_table[9][1] ),
    .A2(\dmmu1.page_table[10][1] ),
    .A3(\dmmu1.page_table[11][1] ),
    .S0(_0891_),
    .S1(_0860_),
    .X(_0935_));
 sky130_fd_sc_hd__a21o_1 _3344_ (.A1(_0872_),
    .A2(_0935_),
    .B1(_0874_),
    .X(_0936_));
 sky130_fd_sc_hd__mux4_1 _3345_ (.A0(\dmmu1.page_table[0][1] ),
    .A1(\dmmu1.page_table[1][1] ),
    .A2(\dmmu1.page_table[2][1] ),
    .A3(\dmmu1.page_table[3][1] ),
    .S0(_0891_),
    .S1(_0860_),
    .X(_0937_));
 sky130_fd_sc_hd__a21o_1 _3346_ (.A1(_0881_),
    .A2(_0937_),
    .B1(_0887_),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_1 _3347_ (.A0(\dmmu1.page_table[6][1] ),
    .A1(\dmmu1.page_table[7][1] ),
    .S(_0858_),
    .X(_0939_));
 sky130_fd_sc_hd__mux2_1 _3348_ (.A0(\dmmu1.page_table[4][1] ),
    .A1(\dmmu1.page_table[5][1] ),
    .S(_0857_),
    .X(_0940_));
 sky130_fd_sc_hd__or2_1 _3349_ (.A(_0863_),
    .B(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__o211a_1 _3350_ (.A1(_0869_),
    .A2(_0939_),
    .B1(_0941_),
    .C1(_0855_),
    .X(_0942_));
 sky130_fd_sc_hd__o22a_1 _3351_ (.A1(_0934_),
    .A2(_0936_),
    .B1(_0938_),
    .B2(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_2 _3352_ (.A0(_0864_),
    .A1(_0943_),
    .S(_0880_),
    .X(_0944_));
 sky130_fd_sc_hd__mux4_1 _3353_ (.A0(\dmmu0.page_table[12][1] ),
    .A1(\dmmu0.page_table[13][1] ),
    .A2(\dmmu0.page_table[14][1] ),
    .A3(\dmmu0.page_table[15][1] ),
    .S0(_0910_),
    .S1(_0913_),
    .X(_0945_));
 sky130_fd_sc_hd__mux4_1 _3354_ (.A0(\dmmu0.page_table[8][1] ),
    .A1(\dmmu0.page_table[9][1] ),
    .A2(\dmmu0.page_table[10][1] ),
    .A3(\dmmu0.page_table[11][1] ),
    .S0(_0910_),
    .S1(_0913_),
    .X(_0946_));
 sky130_fd_sc_hd__mux2_2 _3355_ (.A0(_0945_),
    .A1(_0946_),
    .S(_0918_),
    .X(_0947_));
 sky130_fd_sc_hd__buf_4 _3356_ (.A(_0913_),
    .X(_0948_));
 sky130_fd_sc_hd__mux4_1 _3357_ (.A0(\dmmu0.page_table[4][1] ),
    .A1(\dmmu0.page_table[5][1] ),
    .A2(\dmmu0.page_table[6][1] ),
    .A3(\dmmu0.page_table[7][1] ),
    .S0(_0898_),
    .S1(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__mux2_1 _3358_ (.A0(\dmmu0.page_table[0][1] ),
    .A1(\dmmu0.page_table[1][1] ),
    .S(_0910_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _3359_ (.A0(\dmmu0.page_table[2][1] ),
    .A1(\dmmu0.page_table[3][1] ),
    .S(_0900_),
    .X(_0951_));
 sky130_fd_sc_hd__or2_1 _3360_ (.A(_0909_),
    .B(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__o211a_1 _3361_ (.A1(_0948_),
    .A2(_0950_),
    .B1(_0952_),
    .C1(_0918_),
    .X(_0953_));
 sky130_fd_sc_hd__a211o_1 _3362_ (.A1(_0906_),
    .A2(_0949_),
    .B1(_0953_),
    .C1(_0899_),
    .X(_0954_));
 sky130_fd_sc_hd__o21ai_1 _3363_ (.A1(_0921_),
    .A2(_0947_),
    .B1(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__nand2_1 _3364_ (.A(_0929_),
    .B(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__clkbuf_4 _3365_ (.A(_0927_),
    .X(_0957_));
 sky130_fd_sc_hd__or2_1 _3366_ (.A(_0957_),
    .B(_0928_),
    .X(_0958_));
 sky130_fd_sc_hd__a21oi_1 _3367_ (.A1(_0909_),
    .A2(_0958_),
    .B1(_0819_),
    .Y(_0959_));
 sky130_fd_sc_hd__a22o_2 _3368_ (.A1(_0819_),
    .A2(_0944_),
    .B1(_0956_),
    .B2(_0959_),
    .X(net524));
 sky130_fd_sc_hd__mux4_1 _3369_ (.A0(\dmmu1.page_table[4][2] ),
    .A1(\dmmu1.page_table[5][2] ),
    .A2(\dmmu1.page_table[6][2] ),
    .A3(\dmmu1.page_table[7][2] ),
    .S0(_0892_),
    .S1(_0864_),
    .X(_0960_));
 sky130_fd_sc_hd__mux4_1 _3370_ (.A0(\dmmu1.page_table[12][2] ),
    .A1(\dmmu1.page_table[13][2] ),
    .A2(\dmmu1.page_table[14][2] ),
    .A3(\dmmu1.page_table[15][2] ),
    .S0(_0892_),
    .S1(_0864_),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_1 _3371_ (.A0(_0960_),
    .A1(_0961_),
    .S(_0887_),
    .X(_0962_));
 sky130_fd_sc_hd__o21a_2 _3372_ (.A1(_0893_),
    .A2(_0962_),
    .B1(_0855_),
    .X(_0963_));
 sky130_fd_sc_hd__mux4_1 _3373_ (.A0(\dmmu1.page_table[0][2] ),
    .A1(\dmmu1.page_table[1][2] ),
    .A2(\dmmu1.page_table[2][2] ),
    .A3(\dmmu1.page_table[3][2] ),
    .S0(_0892_),
    .S1(_0864_),
    .X(_0964_));
 sky130_fd_sc_hd__mux4_1 _3374_ (.A0(\dmmu1.page_table[8][2] ),
    .A1(\dmmu1.page_table[9][2] ),
    .A2(\dmmu1.page_table[10][2] ),
    .A3(\dmmu1.page_table[11][2] ),
    .S0(_0892_),
    .S1(_0861_),
    .X(_0965_));
 sky130_fd_sc_hd__mux2_1 _3375_ (.A0(_0964_),
    .A1(_0965_),
    .S(_0887_),
    .X(_0966_));
 sky130_fd_sc_hd__a31o_2 _3376_ (.A1(_0881_),
    .A2(_0880_),
    .A3(_0966_),
    .B1(_0840_),
    .X(_0967_));
 sky130_fd_sc_hd__mux4_1 _3377_ (.A0(\dmmu0.page_table[12][2] ),
    .A1(\dmmu0.page_table[13][2] ),
    .A2(\dmmu0.page_table[14][2] ),
    .A3(\dmmu0.page_table[15][2] ),
    .S0(_0898_),
    .S1(_0948_),
    .X(_0968_));
 sky130_fd_sc_hd__and2_1 _3378_ (.A(_0899_),
    .B(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__mux4_1 _3379_ (.A0(\dmmu0.page_table[4][2] ),
    .A1(\dmmu0.page_table[5][2] ),
    .A2(\dmmu0.page_table[6][2] ),
    .A3(\dmmu0.page_table[7][2] ),
    .S0(_0898_),
    .S1(_0948_),
    .X(_0970_));
 sky130_fd_sc_hd__and2_1 _3380_ (.A(_0921_),
    .B(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__o31a_1 _3381_ (.A1(_0958_),
    .A2(_0969_),
    .A3(_0971_),
    .B1(_0906_),
    .X(_0972_));
 sky130_fd_sc_hd__mux4_1 _3382_ (.A0(\dmmu0.page_table[0][2] ),
    .A1(\dmmu0.page_table[1][2] ),
    .A2(\dmmu0.page_table[2][2] ),
    .A3(\dmmu0.page_table[3][2] ),
    .S0(_0898_),
    .S1(_0948_),
    .X(_0973_));
 sky130_fd_sc_hd__mux4_1 _3383_ (.A0(\dmmu0.page_table[8][2] ),
    .A1(\dmmu0.page_table[9][2] ),
    .A2(\dmmu0.page_table[10][2] ),
    .A3(\dmmu0.page_table[11][2] ),
    .S0(_0898_),
    .S1(_0948_),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_1 _3384_ (.A0(_0973_),
    .A1(_0974_),
    .S(_0899_),
    .X(_0975_));
 sky130_fd_sc_hd__a31o_1 _3385_ (.A1(_0918_),
    .A2(_0929_),
    .A3(_0975_),
    .B1(_0835_),
    .X(_0976_));
 sky130_fd_sc_hd__o22a_2 _3386_ (.A1(_0963_),
    .A2(_0967_),
    .B1(_0972_),
    .B2(_0976_),
    .X(net525));
 sky130_fd_sc_hd__mux4_1 _3387_ (.A0(\dmmu1.page_table[8][3] ),
    .A1(\dmmu1.page_table[9][3] ),
    .A2(\dmmu1.page_table[10][3] ),
    .A3(\dmmu1.page_table[11][3] ),
    .S0(_0892_),
    .S1(_0864_),
    .X(_0977_));
 sky130_fd_sc_hd__mux4_1 _3388_ (.A0(\dmmu1.page_table[12][3] ),
    .A1(\dmmu1.page_table[13][3] ),
    .A2(\dmmu1.page_table[14][3] ),
    .A3(\dmmu1.page_table[15][3] ),
    .S0(_0892_),
    .S1(_0864_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _3389_ (.A0(_0977_),
    .A1(_0978_),
    .S(_0855_),
    .X(_0979_));
 sky130_fd_sc_hd__o21a_2 _3390_ (.A1(_0893_),
    .A2(_0979_),
    .B1(_0887_),
    .X(_0980_));
 sky130_fd_sc_hd__mux4_1 _3391_ (.A0(\dmmu1.page_table[0][3] ),
    .A1(\dmmu1.page_table[1][3] ),
    .A2(\dmmu1.page_table[2][3] ),
    .A3(\dmmu1.page_table[3][3] ),
    .S0(_0892_),
    .S1(_0864_),
    .X(_0981_));
 sky130_fd_sc_hd__mux4_1 _3392_ (.A0(\dmmu1.page_table[4][3] ),
    .A1(\dmmu1.page_table[5][3] ),
    .A2(\dmmu1.page_table[6][3] ),
    .A3(\dmmu1.page_table[7][3] ),
    .S0(_0858_),
    .S1(_0861_),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _3393_ (.A0(_0981_),
    .A1(_0982_),
    .S(_0855_),
    .X(_0983_));
 sky130_fd_sc_hd__a31o_2 _3394_ (.A1(_0874_),
    .A2(_0880_),
    .A3(_0983_),
    .B1(_0840_),
    .X(_0984_));
 sky130_fd_sc_hd__mux4_1 _3395_ (.A0(\dmmu0.page_table[0][3] ),
    .A1(\dmmu0.page_table[1][3] ),
    .A2(\dmmu0.page_table[2][3] ),
    .A3(\dmmu0.page_table[3][3] ),
    .S0(_0898_),
    .S1(_0913_),
    .X(_0985_));
 sky130_fd_sc_hd__mux4_1 _3396_ (.A0(\dmmu0.page_table[4][3] ),
    .A1(\dmmu0.page_table[5][3] ),
    .A2(\dmmu0.page_table[6][3] ),
    .A3(\dmmu0.page_table[7][3] ),
    .S0(_0910_),
    .S1(_0913_),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_1 _3397_ (.A0(_0985_),
    .A1(_0986_),
    .S(_0906_),
    .X(_0987_));
 sky130_fd_sc_hd__a31o_1 _3398_ (.A1(_0921_),
    .A2(_0929_),
    .A3(_0987_),
    .B1(_0835_),
    .X(_0988_));
 sky130_fd_sc_hd__mux4_1 _3399_ (.A0(\dmmu0.page_table[8][3] ),
    .A1(\dmmu0.page_table[9][3] ),
    .A2(\dmmu0.page_table[10][3] ),
    .A3(\dmmu0.page_table[11][3] ),
    .S0(_0898_),
    .S1(_0948_),
    .X(_0989_));
 sky130_fd_sc_hd__mux4_1 _3400_ (.A0(\dmmu0.page_table[12][3] ),
    .A1(\dmmu0.page_table[13][3] ),
    .A2(\dmmu0.page_table[14][3] ),
    .A3(\dmmu0.page_table[15][3] ),
    .S0(_0898_),
    .S1(_0948_),
    .X(_0990_));
 sky130_fd_sc_hd__mux2_1 _3401_ (.A0(_0989_),
    .A1(_0990_),
    .S(_0906_),
    .X(_0991_));
 sky130_fd_sc_hd__o21a_1 _3402_ (.A1(_0958_),
    .A2(_0991_),
    .B1(_0899_),
    .X(_0992_));
 sky130_fd_sc_hd__o22a_4 _3403_ (.A1(_0980_),
    .A2(_0984_),
    .B1(_0988_),
    .B2(_0992_),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_4 _3404_ (.A(_0839_),
    .X(_0993_));
 sky130_fd_sc_hd__inv_2 _3405_ (.A(net158),
    .Y(_0994_));
 sky130_fd_sc_hd__and2_1 _3406_ (.A(net106),
    .B(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__nor3_1 _3407_ (.A(_0994_),
    .B(_0876_),
    .C(_0877_),
    .Y(_0996_));
 sky130_fd_sc_hd__mux4_1 _3408_ (.A0(\dmmu1.page_table[12][4] ),
    .A1(\dmmu1.page_table[13][4] ),
    .A2(\dmmu1.page_table[14][4] ),
    .A3(\dmmu1.page_table[15][4] ),
    .S0(_0891_),
    .S1(_0860_),
    .X(_0997_));
 sky130_fd_sc_hd__or2_1 _3409_ (.A(_0872_),
    .B(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__mux4_1 _3410_ (.A0(\dmmu1.page_table[8][4] ),
    .A1(\dmmu1.page_table[9][4] ),
    .A2(\dmmu1.page_table[10][4] ),
    .A3(\dmmu1.page_table[11][4] ),
    .S0(_0891_),
    .S1(_0860_),
    .X(_0999_));
 sky130_fd_sc_hd__or2_1 _3411_ (.A(_0855_),
    .B(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__mux4_1 _3412_ (.A0(\dmmu1.page_table[0][4] ),
    .A1(\dmmu1.page_table[1][4] ),
    .A2(\dmmu1.page_table[2][4] ),
    .A3(\dmmu1.page_table[3][4] ),
    .S0(_0865_),
    .S1(_0863_),
    .X(_1001_));
 sky130_fd_sc_hd__or2_1 _3413_ (.A(_0855_),
    .B(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__mux4_1 _3414_ (.A0(\dmmu1.page_table[4][4] ),
    .A1(\dmmu1.page_table[5][4] ),
    .A2(\dmmu1.page_table[6][4] ),
    .A3(\dmmu1.page_table[7][4] ),
    .S0(_0865_),
    .S1(_0863_),
    .X(_1003_));
 sky130_fd_sc_hd__o21a_1 _3415_ (.A1(_0881_),
    .A2(_1003_),
    .B1(_0874_),
    .X(_1004_));
 sky130_fd_sc_hd__a32o_2 _3416_ (.A1(_0887_),
    .A2(_0998_),
    .A3(_1000_),
    .B1(_1002_),
    .B2(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__o21a_2 _3417_ (.A1(_0995_),
    .A2(_0996_),
    .B1(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__and2b_2 _3418_ (.A_N(_0995_),
    .B(net124),
    .X(_1007_));
 sky130_fd_sc_hd__nor2_1 _3419_ (.A(_0924_),
    .B(_0925_),
    .Y(_1008_));
 sky130_fd_sc_hd__and2b_1 _3420_ (.A_N(net53),
    .B(net1),
    .X(_1009_));
 sky130_fd_sc_hd__a21o_1 _3421_ (.A1(net53),
    .A2(_1008_),
    .B1(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__mux4_1 _3422_ (.A0(\dmmu0.page_table[8][4] ),
    .A1(\dmmu0.page_table[9][4] ),
    .A2(\dmmu0.page_table[10][4] ),
    .A3(\dmmu0.page_table[11][4] ),
    .S0(_0897_),
    .S1(_0913_),
    .X(_1011_));
 sky130_fd_sc_hd__or2_1 _3423_ (.A(_0906_),
    .B(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__mux4_1 _3424_ (.A0(\dmmu0.page_table[12][4] ),
    .A1(\dmmu0.page_table[13][4] ),
    .A2(\dmmu0.page_table[14][4] ),
    .A3(\dmmu0.page_table[15][4] ),
    .S0(_0897_),
    .S1(_0913_),
    .X(_1013_));
 sky130_fd_sc_hd__o21a_1 _3425_ (.A1(_0918_),
    .A2(_1013_),
    .B1(_0899_),
    .X(_1014_));
 sky130_fd_sc_hd__mux4_1 _3426_ (.A0(\dmmu0.page_table[0][4] ),
    .A1(\dmmu0.page_table[1][4] ),
    .A2(\dmmu0.page_table[2][4] ),
    .A3(\dmmu0.page_table[3][4] ),
    .S0(_0897_),
    .S1(_0902_),
    .X(_1015_));
 sky130_fd_sc_hd__mux4_1 _3427_ (.A0(\dmmu0.page_table[4][4] ),
    .A1(\dmmu0.page_table[5][4] ),
    .A2(\dmmu0.page_table[6][4] ),
    .A3(\dmmu0.page_table[7][4] ),
    .S0(_0897_),
    .S1(_0902_),
    .X(_1016_));
 sky130_fd_sc_hd__mux2_1 _3428_ (.A0(_1015_),
    .A1(_1016_),
    .S(_0906_),
    .X(_1017_));
 sky130_fd_sc_hd__a22o_1 _3429_ (.A1(_1012_),
    .A2(_1014_),
    .B1(_1017_),
    .B2(_0921_),
    .X(_1018_));
 sky130_fd_sc_hd__and2b_1 _3430_ (.A_N(_1009_),
    .B(net19),
    .X(_1019_));
 sky130_fd_sc_hd__a211o_1 _3431_ (.A1(_1010_),
    .A2(_1018_),
    .B1(_1019_),
    .C1(_0835_),
    .X(_1020_));
 sky130_fd_sc_hd__o31a_4 _3432_ (.A1(_0993_),
    .A2(_1006_),
    .A3(_1007_),
    .B1(_1020_),
    .X(net527));
 sky130_fd_sc_hd__mux4_1 _3433_ (.A0(\dmmu1.page_table[0][5] ),
    .A1(\dmmu1.page_table[1][5] ),
    .A2(\dmmu1.page_table[2][5] ),
    .A3(\dmmu1.page_table[3][5] ),
    .S0(_0858_),
    .S1(_0861_),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_1 _3434_ (.A0(\dmmu1.page_table[6][5] ),
    .A1(\dmmu1.page_table[7][5] ),
    .S(_0865_),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_1 _3435_ (.A0(\dmmu1.page_table[4][5] ),
    .A1(\dmmu1.page_table[5][5] ),
    .S(_0857_),
    .X(_1023_));
 sky130_fd_sc_hd__or2_1 _3436_ (.A(_0863_),
    .B(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__o211a_1 _3437_ (.A1(_0869_),
    .A2(_1022_),
    .B1(_1024_),
    .C1(_0855_),
    .X(_1025_));
 sky130_fd_sc_hd__a211o_1 _3438_ (.A1(_0881_),
    .A2(_1021_),
    .B1(_1025_),
    .C1(_0887_),
    .X(_1026_));
 sky130_fd_sc_hd__mux4_1 _3439_ (.A0(\dmmu1.page_table[8][5] ),
    .A1(\dmmu1.page_table[9][5] ),
    .A2(\dmmu1.page_table[10][5] ),
    .A3(\dmmu1.page_table[11][5] ),
    .S0(_0892_),
    .S1(_0864_),
    .X(_1027_));
 sky130_fd_sc_hd__mux2_1 _3440_ (.A0(\dmmu1.page_table[14][5] ),
    .A1(\dmmu1.page_table[15][5] ),
    .S(_0865_),
    .X(_1028_));
 sky130_fd_sc_hd__mux2_1 _3441_ (.A0(\dmmu1.page_table[12][5] ),
    .A1(\dmmu1.page_table[13][5] ),
    .S(_0857_),
    .X(_1029_));
 sky130_fd_sc_hd__or2_1 _3442_ (.A(_0863_),
    .B(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__o211a_1 _3443_ (.A1(_0869_),
    .A2(_1028_),
    .B1(_1030_),
    .C1(_0855_),
    .X(_1031_));
 sky130_fd_sc_hd__a211o_1 _3444_ (.A1(_0881_),
    .A2(_1027_),
    .B1(_1031_),
    .C1(_0874_),
    .X(_1032_));
 sky130_fd_sc_hd__xor2_1 _3445_ (.A(net150),
    .B(\dmmu1.long_off_reg[0] ),
    .X(_1033_));
 sky130_fd_sc_hd__and2_2 _3446_ (.A(net158),
    .B(_0878_),
    .X(_1034_));
 sky130_fd_sc_hd__a32o_2 _3447_ (.A1(_0880_),
    .A2(_1026_),
    .A3(_1032_),
    .B1(_1033_),
    .B2(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _3448_ (.A0(\dmmu0.page_table[6][5] ),
    .A1(\dmmu0.page_table[7][5] ),
    .S(_0898_),
    .X(_1036_));
 sky130_fd_sc_hd__mux2_1 _3449_ (.A0(\dmmu0.page_table[4][5] ),
    .A1(\dmmu0.page_table[5][5] ),
    .S(_0910_),
    .X(_1037_));
 sky130_fd_sc_hd__or2_1 _3450_ (.A(_0948_),
    .B(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__o211a_1 _3451_ (.A1(_0909_),
    .A2(_1036_),
    .B1(_1038_),
    .C1(_0906_),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _3452_ (.A0(\dmmu0.page_table[0][5] ),
    .A1(\dmmu0.page_table[1][5] ),
    .S(_0910_),
    .X(_1040_));
 sky130_fd_sc_hd__or2_1 _3453_ (.A(_0948_),
    .B(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__mux2_1 _3454_ (.A0(\dmmu0.page_table[2][5] ),
    .A1(\dmmu0.page_table[3][5] ),
    .S(_0910_),
    .X(_1042_));
 sky130_fd_sc_hd__or2_1 _3455_ (.A(_0909_),
    .B(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__a31o_1 _3456_ (.A1(_0918_),
    .A2(_1041_),
    .A3(_1043_),
    .B1(_0899_),
    .X(_1044_));
 sky130_fd_sc_hd__mux2_1 _3457_ (.A0(\dmmu0.page_table[10][5] ),
    .A1(\dmmu0.page_table[11][5] ),
    .S(_0910_),
    .X(_1045_));
 sky130_fd_sc_hd__mux2_1 _3458_ (.A0(\dmmu0.page_table[8][5] ),
    .A1(\dmmu0.page_table[9][5] ),
    .S(_0896_),
    .X(_1046_));
 sky130_fd_sc_hd__or2_1 _3459_ (.A(_0913_),
    .B(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__o211a_1 _3460_ (.A1(_0909_),
    .A2(_1045_),
    .B1(_1047_),
    .C1(_0918_),
    .X(_1048_));
 sky130_fd_sc_hd__mux2_1 _3461_ (.A0(\dmmu0.page_table[14][5] ),
    .A1(\dmmu0.page_table[15][5] ),
    .S(_0910_),
    .X(_1049_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(\dmmu0.page_table[12][5] ),
    .A1(\dmmu0.page_table[13][5] ),
    .S(_0900_),
    .X(_1050_));
 sky130_fd_sc_hd__or2_1 _3463_ (.A(_0913_),
    .B(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__o211a_1 _3464_ (.A1(_0909_),
    .A2(_1049_),
    .B1(_1051_),
    .C1(_0906_),
    .X(_1052_));
 sky130_fd_sc_hd__or3_1 _3465_ (.A(_0921_),
    .B(_1048_),
    .C(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__o211a_1 _3466_ (.A1(_1039_),
    .A2(_1044_),
    .B1(_0929_),
    .C1(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__nand2_1 _3467_ (.A(net45),
    .B(\dmmu0.long_off_reg[0] ),
    .Y(_1055_));
 sky130_fd_sc_hd__or2_1 _3468_ (.A(net45),
    .B(\dmmu0.long_off_reg[0] ),
    .X(_1056_));
 sky130_fd_sc_hd__a31o_1 _3469_ (.A1(_0957_),
    .A2(_1055_),
    .A3(_1056_),
    .B1(_0835_),
    .X(_1057_));
 sky130_fd_sc_hd__o22a_4 _3470_ (.A1(_0993_),
    .A2(_1035_),
    .B1(_1054_),
    .B2(_1057_),
    .X(net528));
 sky130_fd_sc_hd__mux4_1 _3471_ (.A0(\dmmu1.page_table[4][6] ),
    .A1(\dmmu1.page_table[5][6] ),
    .A2(\dmmu1.page_table[6][6] ),
    .A3(\dmmu1.page_table[7][6] ),
    .S0(_0858_),
    .S1(_0861_),
    .X(_1058_));
 sky130_fd_sc_hd__mux4_1 _3472_ (.A0(\dmmu1.page_table[0][6] ),
    .A1(\dmmu1.page_table[1][6] ),
    .A2(\dmmu1.page_table[2][6] ),
    .A3(\dmmu1.page_table[3][6] ),
    .S0(_0858_),
    .S1(_0861_),
    .X(_1059_));
 sky130_fd_sc_hd__mux2_1 _3473_ (.A0(_1058_),
    .A1(_1059_),
    .S(_0881_),
    .X(_1060_));
 sky130_fd_sc_hd__mux4_1 _3474_ (.A0(\dmmu1.page_table[12][6] ),
    .A1(\dmmu1.page_table[13][6] ),
    .A2(\dmmu1.page_table[14][6] ),
    .A3(\dmmu1.page_table[15][6] ),
    .S0(_0858_),
    .S1(_0861_),
    .X(_1061_));
 sky130_fd_sc_hd__mux4_1 _3475_ (.A0(\dmmu1.page_table[8][6] ),
    .A1(\dmmu1.page_table[9][6] ),
    .A2(\dmmu1.page_table[10][6] ),
    .A3(\dmmu1.page_table[11][6] ),
    .S0(_0858_),
    .S1(_0861_),
    .X(_1062_));
 sky130_fd_sc_hd__mux2_1 _3476_ (.A0(_1061_),
    .A1(_1062_),
    .S(_0881_),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_1 _3477_ (.A0(_1060_),
    .A1(_1063_),
    .S(_0887_),
    .X(_1064_));
 sky130_fd_sc_hd__nand2_2 _3478_ (.A(_0880_),
    .B(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__xor2_1 _3479_ (.A(net151),
    .B(\dmmu1.long_off_reg[1] ),
    .X(_1066_));
 sky130_fd_sc_hd__a21oi_1 _3480_ (.A1(net150),
    .A2(\dmmu1.long_off_reg[0] ),
    .B1(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__and3_1 _3481_ (.A(net150),
    .B(\dmmu1.long_off_reg[0] ),
    .C(_1066_),
    .X(_1068_));
 sky130_fd_sc_hd__o31a_2 _3482_ (.A1(_0879_),
    .A2(_1067_),
    .A3(_1068_),
    .B1(_0819_),
    .X(_1069_));
 sky130_fd_sc_hd__mux4_1 _3483_ (.A0(\dmmu0.page_table[4][6] ),
    .A1(\dmmu0.page_table[5][6] ),
    .A2(\dmmu0.page_table[6][6] ),
    .A3(\dmmu0.page_table[7][6] ),
    .S0(_0900_),
    .S1(_0902_),
    .X(_1070_));
 sky130_fd_sc_hd__mux4_1 _3484_ (.A0(\dmmu0.page_table[0][6] ),
    .A1(\dmmu0.page_table[1][6] ),
    .A2(\dmmu0.page_table[2][6] ),
    .A3(\dmmu0.page_table[3][6] ),
    .S0(_0900_),
    .S1(_0912_),
    .X(_1071_));
 sky130_fd_sc_hd__mux2_1 _3485_ (.A0(_1070_),
    .A1(_1071_),
    .S(_0918_),
    .X(_1072_));
 sky130_fd_sc_hd__mux4_1 _3486_ (.A0(\dmmu0.page_table[12][6] ),
    .A1(\dmmu0.page_table[13][6] ),
    .A2(\dmmu0.page_table[14][6] ),
    .A3(\dmmu0.page_table[15][6] ),
    .S0(_0900_),
    .S1(_0912_),
    .X(_1073_));
 sky130_fd_sc_hd__mux4_1 _3487_ (.A0(\dmmu0.page_table[8][6] ),
    .A1(\dmmu0.page_table[9][6] ),
    .A2(\dmmu0.page_table[10][6] ),
    .A3(\dmmu0.page_table[11][6] ),
    .S0(_0900_),
    .S1(_0912_),
    .X(_1074_));
 sky130_fd_sc_hd__mux2_1 _3488_ (.A0(_1073_),
    .A1(_1074_),
    .S(_0917_),
    .X(_1075_));
 sky130_fd_sc_hd__mux2_1 _3489_ (.A0(_1072_),
    .A1(_1075_),
    .S(_0899_),
    .X(_1076_));
 sky130_fd_sc_hd__xor2_1 _3490_ (.A(net46),
    .B(\dmmu0.long_off_reg[1] ),
    .X(_1077_));
 sky130_fd_sc_hd__xnor2_1 _3491_ (.A(_1055_),
    .B(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__a22o_1 _3492_ (.A1(_0929_),
    .A2(_1076_),
    .B1(_1078_),
    .B2(_0957_),
    .X(_1079_));
 sky130_fd_sc_hd__o2bb2a_4 _3493_ (.A1_N(_1065_),
    .A2_N(_1069_),
    .B1(_1079_),
    .B2(_0819_),
    .X(net529));
 sky130_fd_sc_hd__mux4_1 _3494_ (.A0(\dmmu1.page_table[4][7] ),
    .A1(\dmmu1.page_table[5][7] ),
    .A2(\dmmu1.page_table[6][7] ),
    .A3(\dmmu1.page_table[7][7] ),
    .S0(_0892_),
    .S1(_0861_),
    .X(_1080_));
 sky130_fd_sc_hd__mux4_1 _3495_ (.A0(\dmmu1.page_table[0][7] ),
    .A1(\dmmu1.page_table[1][7] ),
    .A2(\dmmu1.page_table[2][7] ),
    .A3(\dmmu1.page_table[3][7] ),
    .S0(_0858_),
    .S1(_0861_),
    .X(_1081_));
 sky130_fd_sc_hd__mux2_1 _3496_ (.A0(_1080_),
    .A1(_1081_),
    .S(_0881_),
    .X(_1082_));
 sky130_fd_sc_hd__mux4_1 _3497_ (.A0(\dmmu1.page_table[12][7] ),
    .A1(\dmmu1.page_table[13][7] ),
    .A2(\dmmu1.page_table[14][7] ),
    .A3(\dmmu1.page_table[15][7] ),
    .S0(_0891_),
    .S1(_0860_),
    .X(_1083_));
 sky130_fd_sc_hd__mux4_1 _3498_ (.A0(\dmmu1.page_table[8][7] ),
    .A1(\dmmu1.page_table[9][7] ),
    .A2(\dmmu1.page_table[10][7] ),
    .A3(\dmmu1.page_table[11][7] ),
    .S0(_0891_),
    .S1(_0860_),
    .X(_1084_));
 sky130_fd_sc_hd__mux2_1 _3499_ (.A0(_1083_),
    .A1(_1084_),
    .S(_0872_),
    .X(_1085_));
 sky130_fd_sc_hd__and2_1 _3500_ (.A(_0887_),
    .B(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__a211o_2 _3501_ (.A1(_0874_),
    .A2(_1082_),
    .B1(_1086_),
    .C1(_1034_),
    .X(_1087_));
 sky130_fd_sc_hd__o21a_2 _3502_ (.A1(net106),
    .A2(net158),
    .B1(_0835_),
    .X(_1088_));
 sky130_fd_sc_hd__nand2_1 _3503_ (.A(net152),
    .B(\dmmu1.long_off_reg[2] ),
    .Y(_1089_));
 sky130_fd_sc_hd__or2_1 _3504_ (.A(net152),
    .B(\dmmu1.long_off_reg[2] ),
    .X(_1090_));
 sky130_fd_sc_hd__and2_1 _3505_ (.A(net151),
    .B(\dmmu1.long_off_reg[1] ),
    .X(_1091_));
 sky130_fd_sc_hd__a31o_1 _3506_ (.A1(net150),
    .A2(\dmmu1.long_off_reg[0] ),
    .A3(_1066_),
    .B1(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__a21oi_1 _3507_ (.A1(_1089_),
    .A2(_1090_),
    .B1(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__and3_1 _3508_ (.A(_1089_),
    .B(_1090_),
    .C(_1092_),
    .X(_1094_));
 sky130_fd_sc_hd__o21ai_2 _3509_ (.A1(_1093_),
    .A2(_1094_),
    .B1(_1034_),
    .Y(_1095_));
 sky130_fd_sc_hd__mux4_1 _3510_ (.A0(\dmmu0.page_table[4][7] ),
    .A1(\dmmu0.page_table[5][7] ),
    .A2(\dmmu0.page_table[6][7] ),
    .A3(\dmmu0.page_table[7][7] ),
    .S0(_0897_),
    .S1(_0902_),
    .X(_1096_));
 sky130_fd_sc_hd__mux4_1 _3511_ (.A0(\dmmu0.page_table[0][7] ),
    .A1(\dmmu0.page_table[1][7] ),
    .A2(\dmmu0.page_table[2][7] ),
    .A3(\dmmu0.page_table[3][7] ),
    .S0(_0897_),
    .S1(_0902_),
    .X(_1097_));
 sky130_fd_sc_hd__mux2_1 _3512_ (.A0(_1096_),
    .A1(_1097_),
    .S(_0918_),
    .X(_1098_));
 sky130_fd_sc_hd__mux4_1 _3513_ (.A0(\dmmu0.page_table[12][7] ),
    .A1(\dmmu0.page_table[13][7] ),
    .A2(\dmmu0.page_table[14][7] ),
    .A3(\dmmu0.page_table[15][7] ),
    .S0(_0896_),
    .S1(_0912_),
    .X(_1099_));
 sky130_fd_sc_hd__mux4_1 _3514_ (.A0(\dmmu0.page_table[8][7] ),
    .A1(\dmmu0.page_table[9][7] ),
    .A2(\dmmu0.page_table[10][7] ),
    .A3(\dmmu0.page_table[11][7] ),
    .S0(_0896_),
    .S1(_0901_),
    .X(_1100_));
 sky130_fd_sc_hd__mux2_1 _3515_ (.A0(_1099_),
    .A1(_1100_),
    .S(_0917_),
    .X(_1101_));
 sky130_fd_sc_hd__and2_1 _3516_ (.A(_0899_),
    .B(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__a211o_1 _3517_ (.A1(_0921_),
    .A2(_1098_),
    .B1(_1102_),
    .C1(_0957_),
    .X(_1103_));
 sky130_fd_sc_hd__nor2_1 _3518_ (.A(_0818_),
    .B(_0928_),
    .Y(_1104_));
 sky130_fd_sc_hd__and2_1 _3519_ (.A(net47),
    .B(\dmmu0.long_off_reg[2] ),
    .X(_1105_));
 sky130_fd_sc_hd__nor2_1 _3520_ (.A(net47),
    .B(\dmmu0.long_off_reg[2] ),
    .Y(_1106_));
 sky130_fd_sc_hd__and2_1 _3521_ (.A(net46),
    .B(\dmmu0.long_off_reg[1] ),
    .X(_1107_));
 sky130_fd_sc_hd__a31oi_2 _3522_ (.A1(net45),
    .A2(\dmmu0.long_off_reg[0] ),
    .A3(_1077_),
    .B1(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__o21a_1 _3523_ (.A1(_1105_),
    .A2(_1106_),
    .B1(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__nor3_1 _3524_ (.A(_1105_),
    .B(_1106_),
    .C(_1108_),
    .Y(_1110_));
 sky130_fd_sc_hd__o21ai_1 _3525_ (.A1(_1109_),
    .A2(_1110_),
    .B1(_0957_),
    .Y(_1111_));
 sky130_fd_sc_hd__and3_1 _3526_ (.A(_1103_),
    .B(_1104_),
    .C(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__a31o_4 _3527_ (.A1(_1087_),
    .A2(_1088_),
    .A3(_1095_),
    .B1(_1112_),
    .X(net530));
 sky130_fd_sc_hd__mux4_1 _3528_ (.A0(\dmmu1.page_table[0][8] ),
    .A1(\dmmu1.page_table[1][8] ),
    .A2(\dmmu1.page_table[2][8] ),
    .A3(\dmmu1.page_table[3][8] ),
    .S0(_0891_),
    .S1(_0860_),
    .X(_1113_));
 sky130_fd_sc_hd__mux4_1 _3529_ (.A0(\dmmu1.page_table[4][8] ),
    .A1(\dmmu1.page_table[5][8] ),
    .A2(\dmmu1.page_table[6][8] ),
    .A3(\dmmu1.page_table[7][8] ),
    .S0(_0891_),
    .S1(_0860_),
    .X(_1114_));
 sky130_fd_sc_hd__mux2_1 _3530_ (.A0(_1113_),
    .A1(_1114_),
    .S(_0854_),
    .X(_1115_));
 sky130_fd_sc_hd__mux2_1 _3531_ (.A0(\dmmu1.page_table[12][8] ),
    .A1(\dmmu1.page_table[13][8] ),
    .S(_0857_),
    .X(_1116_));
 sky130_fd_sc_hd__or2_1 _3532_ (.A(_0863_),
    .B(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__mux2_1 _3533_ (.A0(\dmmu1.page_table[14][8] ),
    .A1(\dmmu1.page_table[15][8] ),
    .S(_0891_),
    .X(_1118_));
 sky130_fd_sc_hd__o21a_1 _3534_ (.A1(_0869_),
    .A2(_1118_),
    .B1(_0854_),
    .X(_1119_));
 sky130_fd_sc_hd__mux4_1 _3535_ (.A0(\dmmu1.page_table[8][8] ),
    .A1(\dmmu1.page_table[9][8] ),
    .A2(\dmmu1.page_table[10][8] ),
    .A3(\dmmu1.page_table[11][8] ),
    .S0(_0865_),
    .S1(_0863_),
    .X(_1120_));
 sky130_fd_sc_hd__a221o_1 _3536_ (.A1(_1117_),
    .A2(_1119_),
    .B1(_1120_),
    .B2(_0881_),
    .C1(_0874_),
    .X(_1121_));
 sky130_fd_sc_hd__o21a_2 _3537_ (.A1(_0887_),
    .A2(_1115_),
    .B1(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__nand2_1 _3538_ (.A(net153),
    .B(\dmmu1.long_off_reg[3] ),
    .Y(_1123_));
 sky130_fd_sc_hd__or2_1 _3539_ (.A(net153),
    .B(\dmmu1.long_off_reg[3] ),
    .X(_1124_));
 sky130_fd_sc_hd__a21bo_1 _3540_ (.A1(_1090_),
    .A2(_1092_),
    .B1_N(_1089_),
    .X(_1125_));
 sky130_fd_sc_hd__a31oi_1 _3541_ (.A1(_1123_),
    .A2(_1124_),
    .A3(_1125_),
    .B1(_0879_),
    .Y(_1126_));
 sky130_fd_sc_hd__a21o_1 _3542_ (.A1(_1123_),
    .A2(_1124_),
    .B1(_1125_),
    .X(_1127_));
 sky130_fd_sc_hd__a22o_1 _3543_ (.A1(_0879_),
    .A2(_1122_),
    .B1(_1126_),
    .B2(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__nand2_1 _3544_ (.A(net48),
    .B(\dmmu0.long_off_reg[3] ),
    .Y(_1129_));
 sky130_fd_sc_hd__or2_1 _3545_ (.A(net48),
    .B(\dmmu0.long_off_reg[3] ),
    .X(_1130_));
 sky130_fd_sc_hd__o21bai_1 _3546_ (.A1(_1106_),
    .A2(_1108_),
    .B1_N(_1105_),
    .Y(_1131_));
 sky130_fd_sc_hd__a21oi_1 _3547_ (.A1(_1129_),
    .A2(_1130_),
    .B1(_1131_),
    .Y(_1132_));
 sky130_fd_sc_hd__and3_1 _3548_ (.A(_1129_),
    .B(_1130_),
    .C(_1131_),
    .X(_1133_));
 sky130_fd_sc_hd__o21ai_1 _3549_ (.A1(_1132_),
    .A2(_1133_),
    .B1(_0957_),
    .Y(_1134_));
 sky130_fd_sc_hd__mux4_1 _3550_ (.A0(\dmmu0.page_table[4][8] ),
    .A1(\dmmu0.page_table[5][8] ),
    .A2(\dmmu0.page_table[6][8] ),
    .A3(\dmmu0.page_table[7][8] ),
    .S0(_0897_),
    .S1(_0902_),
    .X(_1135_));
 sky130_fd_sc_hd__mux4_1 _3551_ (.A0(\dmmu0.page_table[0][8] ),
    .A1(\dmmu0.page_table[1][8] ),
    .A2(\dmmu0.page_table[2][8] ),
    .A3(\dmmu0.page_table[3][8] ),
    .S0(_0897_),
    .S1(_0902_),
    .X(_1136_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(_1135_),
    .A1(_1136_),
    .S(_0918_),
    .X(_1137_));
 sky130_fd_sc_hd__mux4_1 _3553_ (.A0(\dmmu0.page_table[12][8] ),
    .A1(\dmmu0.page_table[13][8] ),
    .A2(\dmmu0.page_table[14][8] ),
    .A3(\dmmu0.page_table[15][8] ),
    .S0(_0896_),
    .S1(_0912_),
    .X(_1138_));
 sky130_fd_sc_hd__mux4_1 _3554_ (.A0(\dmmu0.page_table[8][8] ),
    .A1(\dmmu0.page_table[9][8] ),
    .A2(\dmmu0.page_table[10][8] ),
    .A3(\dmmu0.page_table[11][8] ),
    .S0(_0896_),
    .S1(_0912_),
    .X(_1139_));
 sky130_fd_sc_hd__mux2_2 _3555_ (.A0(_1138_),
    .A1(_1139_),
    .S(_0917_),
    .X(_1140_));
 sky130_fd_sc_hd__and2_1 _3556_ (.A(_0899_),
    .B(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__a211o_1 _3557_ (.A1(_0921_),
    .A2(_1137_),
    .B1(_1141_),
    .C1(_0957_),
    .X(_1142_));
 sky130_fd_sc_hd__and3_1 _3558_ (.A(_1104_),
    .B(_1134_),
    .C(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__a21o_4 _3559_ (.A1(_1088_),
    .A2(_1128_),
    .B1(_1143_),
    .X(net531));
 sky130_fd_sc_hd__mux2_1 _3560_ (.A0(\dmmu1.page_table[14][9] ),
    .A1(\dmmu1.page_table[15][9] ),
    .S(_0856_),
    .X(_1144_));
 sky130_fd_sc_hd__and2_1 _3561_ (.A(_0859_),
    .B(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__buf_4 _3562_ (.A(_0856_),
    .X(_1146_));
 sky130_fd_sc_hd__mux2_1 _3563_ (.A0(\dmmu1.page_table[12][9] ),
    .A1(\dmmu1.page_table[13][9] ),
    .S(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__a21o_1 _3564_ (.A1(_0868_),
    .A2(_1147_),
    .B1(_0872_),
    .X(_1148_));
 sky130_fd_sc_hd__mux2_1 _3565_ (.A0(\dmmu1.page_table[8][9] ),
    .A1(\dmmu1.page_table[9][9] ),
    .S(_0856_),
    .X(_1149_));
 sky130_fd_sc_hd__and2_1 _3566_ (.A(_0868_),
    .B(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__mux2_1 _3567_ (.A0(\dmmu1.page_table[10][9] ),
    .A1(\dmmu1.page_table[11][9] ),
    .S(_1146_),
    .X(_1151_));
 sky130_fd_sc_hd__a21o_1 _3568_ (.A1(_0859_),
    .A2(_1151_),
    .B1(_0854_),
    .X(_1152_));
 sky130_fd_sc_hd__o221a_2 _3569_ (.A1(_1145_),
    .A2(_1148_),
    .B1(_1150_),
    .B2(_1152_),
    .C1(net123),
    .X(_1153_));
 sky130_fd_sc_hd__mux2_1 _3570_ (.A0(\dmmu1.page_table[4][9] ),
    .A1(\dmmu1.page_table[5][9] ),
    .S(_1146_),
    .X(_1154_));
 sky130_fd_sc_hd__and2_1 _3571_ (.A(_0869_),
    .B(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _3572_ (.A0(\dmmu1.page_table[6][9] ),
    .A1(\dmmu1.page_table[7][9] ),
    .S(_1146_),
    .X(_1156_));
 sky130_fd_sc_hd__a21o_1 _3573_ (.A1(_0859_),
    .A2(_1156_),
    .B1(_0872_),
    .X(_1157_));
 sky130_fd_sc_hd__mux2_1 _3574_ (.A0(\dmmu1.page_table[2][9] ),
    .A1(\dmmu1.page_table[3][9] ),
    .S(_0857_),
    .X(_1158_));
 sky130_fd_sc_hd__mux2_1 _3575_ (.A0(\dmmu1.page_table[0][9] ),
    .A1(\dmmu1.page_table[1][9] ),
    .S(_0856_),
    .X(_1159_));
 sky130_fd_sc_hd__a21o_1 _3576_ (.A1(_0868_),
    .A2(_1159_),
    .B1(_0854_),
    .X(_1160_));
 sky130_fd_sc_hd__a21o_1 _3577_ (.A1(_0859_),
    .A2(_1158_),
    .B1(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__o211a_2 _3578_ (.A1(_1155_),
    .A2(_1157_),
    .B1(_0874_),
    .C1(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__nand2_1 _3579_ (.A(net154),
    .B(\dmmu1.long_off_reg[4] ),
    .Y(_1163_));
 sky130_fd_sc_hd__or2_1 _3580_ (.A(net154),
    .B(\dmmu1.long_off_reg[4] ),
    .X(_1164_));
 sky130_fd_sc_hd__nand2_1 _3581_ (.A(_1163_),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__a21bo_1 _3582_ (.A1(_1124_),
    .A2(_1125_),
    .B1_N(_1123_),
    .X(_1166_));
 sky130_fd_sc_hd__xnor2_1 _3583_ (.A(_1165_),
    .B(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__o32a_2 _3584_ (.A1(_0893_),
    .A2(_1153_),
    .A3(_1162_),
    .B1(_1167_),
    .B2(_0879_),
    .X(_1168_));
 sky130_fd_sc_hd__buf_6 _3585_ (.A(net15),
    .X(_1169_));
 sky130_fd_sc_hd__mux2_1 _3586_ (.A0(\dmmu0.page_table[8][9] ),
    .A1(\dmmu0.page_table[9][9] ),
    .S(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__nand2_1 _3587_ (.A(_0909_),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__mux2_1 _3588_ (.A0(\dmmu0.page_table[10][9] ),
    .A1(\dmmu0.page_table[11][9] ),
    .S(_1169_),
    .X(_1172_));
 sky130_fd_sc_hd__a21oi_1 _3589_ (.A1(_0901_),
    .A2(_1172_),
    .B1(_0905_),
    .Y(_1173_));
 sky130_fd_sc_hd__mux2_1 _3590_ (.A0(\dmmu0.page_table[14][9] ),
    .A1(\dmmu0.page_table[15][9] ),
    .S(_1169_),
    .X(_1174_));
 sky130_fd_sc_hd__nand2_1 _3591_ (.A(_0912_),
    .B(_1174_),
    .Y(_1175_));
 sky130_fd_sc_hd__mux2_1 _3592_ (.A0(\dmmu0.page_table[12][9] ),
    .A1(\dmmu0.page_table[13][9] ),
    .S(_1169_),
    .X(_1176_));
 sky130_fd_sc_hd__a21oi_1 _3593_ (.A1(_0908_),
    .A2(_1176_),
    .B1(_0917_),
    .Y(_1177_));
 sky130_fd_sc_hd__a221o_1 _3594_ (.A1(_1171_),
    .A2(_1173_),
    .B1(_1175_),
    .B2(_1177_),
    .C1(_0921_),
    .X(_1178_));
 sky130_fd_sc_hd__mux2_1 _3595_ (.A0(\dmmu0.page_table[4][9] ),
    .A1(\dmmu0.page_table[5][9] ),
    .S(_1169_),
    .X(_1179_));
 sky130_fd_sc_hd__nand2_1 _3596_ (.A(_0908_),
    .B(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__mux2_1 _3597_ (.A0(\dmmu0.page_table[6][9] ),
    .A1(\dmmu0.page_table[7][9] ),
    .S(_1169_),
    .X(_1181_));
 sky130_fd_sc_hd__nand2_1 _3598_ (.A(_0912_),
    .B(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__mux2_1 _3599_ (.A0(\dmmu0.page_table[2][9] ),
    .A1(\dmmu0.page_table[3][9] ),
    .S(_1169_),
    .X(_1183_));
 sky130_fd_sc_hd__mux2_1 _3600_ (.A0(\dmmu0.page_table[0][9] ),
    .A1(\dmmu0.page_table[1][9] ),
    .S(_0895_),
    .X(_1184_));
 sky130_fd_sc_hd__a21o_1 _3601_ (.A1(_0908_),
    .A2(_1184_),
    .B1(_0905_),
    .X(_1185_));
 sky130_fd_sc_hd__a21oi_1 _3602_ (.A1(_0912_),
    .A2(_1183_),
    .B1(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__a311o_1 _3603_ (.A1(_0905_),
    .A2(_1180_),
    .A3(_1182_),
    .B1(net18),
    .C1(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__nand2_1 _3604_ (.A(net49),
    .B(\dmmu0.long_off_reg[4] ),
    .Y(_1188_));
 sky130_fd_sc_hd__or2_1 _3605_ (.A(net49),
    .B(\dmmu0.long_off_reg[4] ),
    .X(_1189_));
 sky130_fd_sc_hd__nand2_1 _3606_ (.A(_1188_),
    .B(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__a21bo_1 _3607_ (.A1(_1130_),
    .A2(_1131_),
    .B1_N(_1129_),
    .X(_1191_));
 sky130_fd_sc_hd__xor2_1 _3608_ (.A(_1190_),
    .B(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__a32o_1 _3609_ (.A1(_0929_),
    .A2(_1178_),
    .A3(_1187_),
    .B1(_1192_),
    .B2(_0957_),
    .X(_1193_));
 sky130_fd_sc_hd__nand2_1 _3610_ (.A(_0838_),
    .B(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__o21a_4 _3611_ (.A1(_0993_),
    .A2(_1168_),
    .B1(_1194_),
    .X(net533));
 sky130_fd_sc_hd__mux4_1 _3612_ (.A0(\dmmu1.page_table[0][10] ),
    .A1(\dmmu1.page_table[1][10] ),
    .A2(\dmmu1.page_table[2][10] ),
    .A3(\dmmu1.page_table[3][10] ),
    .S0(net120),
    .S1(net121),
    .X(_1195_));
 sky130_fd_sc_hd__mux4_1 _3613_ (.A0(\dmmu1.page_table[4][10] ),
    .A1(\dmmu1.page_table[5][10] ),
    .A2(\dmmu1.page_table[6][10] ),
    .A3(\dmmu1.page_table[7][10] ),
    .S0(net120),
    .S1(net121),
    .X(_1196_));
 sky130_fd_sc_hd__mux2_1 _3614_ (.A0(_1195_),
    .A1(_1196_),
    .S(net122),
    .X(_1197_));
 sky130_fd_sc_hd__mux4_1 _3615_ (.A0(\dmmu1.page_table[8][10] ),
    .A1(\dmmu1.page_table[9][10] ),
    .A2(\dmmu1.page_table[10][10] ),
    .A3(\dmmu1.page_table[11][10] ),
    .S0(net120),
    .S1(net121),
    .X(_1198_));
 sky130_fd_sc_hd__mux2_1 _3616_ (.A0(\dmmu1.page_table[12][10] ),
    .A1(\dmmu1.page_table[13][10] ),
    .S(net120),
    .X(_1199_));
 sky130_fd_sc_hd__or2_1 _3617_ (.A(net121),
    .B(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__mux2_1 _3618_ (.A0(\dmmu1.page_table[14][10] ),
    .A1(\dmmu1.page_table[15][10] ),
    .S(net120),
    .X(_1201_));
 sky130_fd_sc_hd__o21a_1 _3619_ (.A1(_0868_),
    .A2(_1201_),
    .B1(net122),
    .X(_1202_));
 sky130_fd_sc_hd__a221o_1 _3620_ (.A1(_0871_),
    .A2(_1198_),
    .B1(_1200_),
    .B2(_1202_),
    .C1(_0874_),
    .X(_1203_));
 sky130_fd_sc_hd__o21a_2 _3621_ (.A1(net123),
    .A2(_1197_),
    .B1(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__nand2_1 _3622_ (.A(net155),
    .B(\dmmu1.long_off_reg[5] ),
    .Y(_1205_));
 sky130_fd_sc_hd__or2_1 _3623_ (.A(net155),
    .B(\dmmu1.long_off_reg[5] ),
    .X(_1206_));
 sky130_fd_sc_hd__nand2_1 _3624_ (.A(_1205_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__a21boi_1 _3625_ (.A1(_1164_),
    .A2(_1166_),
    .B1_N(_1163_),
    .Y(_1208_));
 sky130_fd_sc_hd__xor2_1 _3626_ (.A(_1207_),
    .B(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__mux2_1 _3627_ (.A0(_1204_),
    .A1(_1209_),
    .S(_0878_),
    .X(_1210_));
 sky130_fd_sc_hd__a22o_2 _3628_ (.A1(_0995_),
    .A2(_1204_),
    .B1(_1210_),
    .B2(net158),
    .X(_1211_));
 sky130_fd_sc_hd__mux2_1 _3629_ (.A0(\dmmu0.page_table[12][10] ),
    .A1(\dmmu0.page_table[13][10] ),
    .S(_0895_),
    .X(_1212_));
 sky130_fd_sc_hd__mux2_1 _3630_ (.A0(\dmmu0.page_table[14][10] ),
    .A1(\dmmu0.page_table[15][10] ),
    .S(net15),
    .X(_1213_));
 sky130_fd_sc_hd__or2_1 _3631_ (.A(_0908_),
    .B(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__o211a_1 _3632_ (.A1(_0901_),
    .A2(_1212_),
    .B1(_1214_),
    .C1(_0905_),
    .X(_1215_));
 sky130_fd_sc_hd__mux4_1 _3633_ (.A0(\dmmu0.page_table[8][10] ),
    .A1(\dmmu0.page_table[9][10] ),
    .A2(\dmmu0.page_table[10][10] ),
    .A3(\dmmu0.page_table[11][10] ),
    .S0(_0895_),
    .S1(net16),
    .X(_1216_));
 sky130_fd_sc_hd__a21o_1 _3634_ (.A1(_0917_),
    .A2(_1216_),
    .B1(_0920_),
    .X(_1217_));
 sky130_fd_sc_hd__mux4_1 _3635_ (.A0(\dmmu0.page_table[0][10] ),
    .A1(\dmmu0.page_table[1][10] ),
    .A2(\dmmu0.page_table[2][10] ),
    .A3(\dmmu0.page_table[3][10] ),
    .S0(_0895_),
    .S1(net16),
    .X(_1218_));
 sky130_fd_sc_hd__mux4_1 _3636_ (.A0(\dmmu0.page_table[4][10] ),
    .A1(\dmmu0.page_table[5][10] ),
    .A2(\dmmu0.page_table[6][10] ),
    .A3(\dmmu0.page_table[7][10] ),
    .S0(net15),
    .S1(net16),
    .X(_1219_));
 sky130_fd_sc_hd__mux2_1 _3637_ (.A0(_1218_),
    .A1(_1219_),
    .S(net17),
    .X(_1220_));
 sky130_fd_sc_hd__o22a_1 _3638_ (.A1(_1215_),
    .A2(_1217_),
    .B1(_1220_),
    .B2(net18),
    .X(_1221_));
 sky130_fd_sc_hd__nand2_1 _3639_ (.A(net50),
    .B(\dmmu0.long_off_reg[5] ),
    .Y(_1222_));
 sky130_fd_sc_hd__or2_1 _3640_ (.A(net50),
    .B(\dmmu0.long_off_reg[5] ),
    .X(_1223_));
 sky130_fd_sc_hd__nand2_1 _3641_ (.A(_1222_),
    .B(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__a21bo_1 _3642_ (.A1(_1189_),
    .A2(_1191_),
    .B1_N(_1188_),
    .X(_1225_));
 sky130_fd_sc_hd__xnor2_1 _3643_ (.A(_1224_),
    .B(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__mux2_1 _3644_ (.A0(_1221_),
    .A1(_1226_),
    .S(_0926_),
    .X(_1227_));
 sky130_fd_sc_hd__a22o_1 _3645_ (.A1(_1009_),
    .A2(_1221_),
    .B1(_1227_),
    .B2(net53),
    .X(_1228_));
 sky130_fd_sc_hd__mux2_4 _3646_ (.A0(_1211_),
    .A1(_1228_),
    .S(_0847_),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _3647_ (.A(_1229_),
    .X(net534));
 sky130_fd_sc_hd__mux2_1 _3648_ (.A0(\dmmu0.page_table[2][11] ),
    .A1(\dmmu0.page_table[3][11] ),
    .S(_1169_),
    .X(_1230_));
 sky130_fd_sc_hd__mux2_1 _3649_ (.A0(\dmmu0.page_table[0][11] ),
    .A1(\dmmu0.page_table[1][11] ),
    .S(_0895_),
    .X(_1231_));
 sky130_fd_sc_hd__or2_1 _3650_ (.A(_0901_),
    .B(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__o211a_1 _3651_ (.A1(_0908_),
    .A2(_1230_),
    .B1(_1232_),
    .C1(_0917_),
    .X(_1233_));
 sky130_fd_sc_hd__mux2_1 _3652_ (.A0(\dmmu0.page_table[6][11] ),
    .A1(\dmmu0.page_table[7][11] ),
    .S(_0896_),
    .X(_1234_));
 sky130_fd_sc_hd__mux2_1 _3653_ (.A0(\dmmu0.page_table[4][11] ),
    .A1(\dmmu0.page_table[5][11] ),
    .S(_0895_),
    .X(_1235_));
 sky130_fd_sc_hd__or2_1 _3654_ (.A(_0901_),
    .B(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__o211a_1 _3655_ (.A1(_0908_),
    .A2(_1234_),
    .B1(_1236_),
    .C1(_0905_),
    .X(_1237_));
 sky130_fd_sc_hd__or3_1 _3656_ (.A(net18),
    .B(_1233_),
    .C(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__mux2_1 _3657_ (.A0(\dmmu0.page_table[10][11] ),
    .A1(\dmmu0.page_table[11][11] ),
    .S(_0896_),
    .X(_1239_));
 sky130_fd_sc_hd__mux2_1 _3658_ (.A0(\dmmu0.page_table[8][11] ),
    .A1(\dmmu0.page_table[9][11] ),
    .S(_0895_),
    .X(_1240_));
 sky130_fd_sc_hd__or2_1 _3659_ (.A(_0901_),
    .B(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__o211a_1 _3660_ (.A1(_0909_),
    .A2(_1239_),
    .B1(_1241_),
    .C1(_0917_),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _3661_ (.A0(\dmmu0.page_table[14][11] ),
    .A1(\dmmu0.page_table[15][11] ),
    .S(_0896_),
    .X(_1243_));
 sky130_fd_sc_hd__mux2_1 _3662_ (.A0(\dmmu0.page_table[12][11] ),
    .A1(\dmmu0.page_table[13][11] ),
    .S(_1169_),
    .X(_1244_));
 sky130_fd_sc_hd__or2_1 _3663_ (.A(_0901_),
    .B(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__o211a_1 _3664_ (.A1(_0909_),
    .A2(_1243_),
    .B1(_1245_),
    .C1(_0905_),
    .X(_1246_));
 sky130_fd_sc_hd__o31a_1 _3665_ (.A1(_0921_),
    .A2(_1242_),
    .A3(_1246_),
    .B1(_0929_),
    .X(_1247_));
 sky130_fd_sc_hd__inv_2 _3666_ (.A(_1222_),
    .Y(_1248_));
 sky130_fd_sc_hd__a21oi_1 _3667_ (.A1(_1223_),
    .A2(_1225_),
    .B1(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__nor2_1 _3668_ (.A(net51),
    .B(\dmmu0.long_off_reg[6] ),
    .Y(_1250_));
 sky130_fd_sc_hd__and2_1 _3669_ (.A(net51),
    .B(\dmmu0.long_off_reg[6] ),
    .X(_1251_));
 sky130_fd_sc_hd__nor2_1 _3670_ (.A(_1250_),
    .B(_1251_),
    .Y(_1252_));
 sky130_fd_sc_hd__xnor2_1 _3671_ (.A(_1249_),
    .B(_1252_),
    .Y(_1253_));
 sky130_fd_sc_hd__a22o_1 _3672_ (.A1(_1238_),
    .A2(_1247_),
    .B1(_1253_),
    .B2(_0957_),
    .X(_1254_));
 sky130_fd_sc_hd__o21ai_1 _3673_ (.A1(_1207_),
    .A2(_1208_),
    .B1(_1205_),
    .Y(_1255_));
 sky130_fd_sc_hd__or2_1 _3674_ (.A(net156),
    .B(\dmmu1.long_off_reg[6] ),
    .X(_1256_));
 sky130_fd_sc_hd__nand2_1 _3675_ (.A(net156),
    .B(\dmmu1.long_off_reg[6] ),
    .Y(_1257_));
 sky130_fd_sc_hd__and3_1 _3676_ (.A(_1255_),
    .B(_1256_),
    .C(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__a21oi_1 _3677_ (.A1(_1256_),
    .A2(_1257_),
    .B1(_1255_),
    .Y(_1259_));
 sky130_fd_sc_hd__mux2_1 _3678_ (.A0(\dmmu1.page_table[8][11] ),
    .A1(\dmmu1.page_table[9][11] ),
    .S(_1146_),
    .X(_1260_));
 sky130_fd_sc_hd__nor2_1 _3679_ (.A(_0859_),
    .B(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__mux2_1 _3680_ (.A0(\dmmu1.page_table[10][11] ),
    .A1(\dmmu1.page_table[11][11] ),
    .S(_0856_),
    .X(_1262_));
 sky130_fd_sc_hd__o21ai_1 _3681_ (.A1(_0868_),
    .A2(_1262_),
    .B1(_0872_),
    .Y(_1263_));
 sky130_fd_sc_hd__mux2_1 _3682_ (.A0(\dmmu1.page_table[14][11] ),
    .A1(\dmmu1.page_table[15][11] ),
    .S(_1146_),
    .X(_1264_));
 sky130_fd_sc_hd__nor2_1 _3683_ (.A(_0869_),
    .B(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__mux2_1 _3684_ (.A0(\dmmu1.page_table[12][11] ),
    .A1(\dmmu1.page_table[13][11] ),
    .S(_1146_),
    .X(_1266_));
 sky130_fd_sc_hd__o21ai_1 _3685_ (.A1(_0859_),
    .A2(_1266_),
    .B1(_0854_),
    .Y(_1267_));
 sky130_fd_sc_hd__o221a_2 _3686_ (.A1(_1261_),
    .A2(_1263_),
    .B1(_1265_),
    .B2(_1267_),
    .C1(net123),
    .X(_1268_));
 sky130_fd_sc_hd__mux2_1 _3687_ (.A0(\dmmu1.page_table[0][11] ),
    .A1(\dmmu1.page_table[1][11] ),
    .S(_0856_),
    .X(_1269_));
 sky130_fd_sc_hd__or2_1 _3688_ (.A(_0859_),
    .B(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_1 _3689_ (.A0(\dmmu1.page_table[2][11] ),
    .A1(\dmmu1.page_table[3][11] ),
    .S(_0856_),
    .X(_1271_));
 sky130_fd_sc_hd__or2_1 _3690_ (.A(_0868_),
    .B(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__mux2_1 _3691_ (.A0(\dmmu1.page_table[6][11] ),
    .A1(\dmmu1.page_table[7][11] ),
    .S(_0856_),
    .X(_1273_));
 sky130_fd_sc_hd__mux2_1 _3692_ (.A0(\dmmu1.page_table[4][11] ),
    .A1(\dmmu1.page_table[5][11] ),
    .S(net120),
    .X(_1274_));
 sky130_fd_sc_hd__or2_1 _3693_ (.A(net121),
    .B(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__o211a_1 _3694_ (.A1(_0868_),
    .A2(_1273_),
    .B1(_1275_),
    .C1(_0854_),
    .X(_1276_));
 sky130_fd_sc_hd__a311o_2 _3695_ (.A1(_0872_),
    .A2(_1270_),
    .A3(_1272_),
    .B1(_1276_),
    .C1(net123),
    .X(_1277_));
 sky130_fd_sc_hd__or3b_1 _3696_ (.A(_0893_),
    .B(_1268_),
    .C_N(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__o31ai_4 _3697_ (.A1(_0879_),
    .A2(_1258_),
    .A3(_1259_),
    .B1(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__mux2_4 _3698_ (.A0(_1254_),
    .A1(_1279_),
    .S(_0835_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _3699_ (.A(_1280_),
    .X(net535));
 sky130_fd_sc_hd__xnor2_1 _3700_ (.A(net52),
    .B(\dmmu0.long_off_reg[7] ),
    .Y(_1281_));
 sky130_fd_sc_hd__a211oi_1 _3701_ (.A1(_1223_),
    .A2(_1225_),
    .B1(_1251_),
    .C1(_1248_),
    .Y(_1282_));
 sky130_fd_sc_hd__or3_1 _3702_ (.A(_1250_),
    .B(_1281_),
    .C(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__o21ai_1 _3703_ (.A1(_1250_),
    .A2(_1282_),
    .B1(_1281_),
    .Y(_1284_));
 sky130_fd_sc_hd__mux4_1 _3704_ (.A0(\dmmu0.page_table[8][12] ),
    .A1(\dmmu0.page_table[9][12] ),
    .A2(\dmmu0.page_table[10][12] ),
    .A3(\dmmu0.page_table[11][12] ),
    .S0(net15),
    .S1(net16),
    .X(_1285_));
 sky130_fd_sc_hd__inv_2 _3705_ (.A(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__mux2_1 _3706_ (.A0(\dmmu0.page_table[12][12] ),
    .A1(\dmmu0.page_table[13][12] ),
    .S(_1169_),
    .X(_1287_));
 sky130_fd_sc_hd__nor2_1 _3707_ (.A(_0901_),
    .B(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hd__mux2_1 _3708_ (.A0(\dmmu0.page_table[14][12] ),
    .A1(\dmmu0.page_table[15][12] ),
    .S(_0895_),
    .X(_1289_));
 sky130_fd_sc_hd__o21ai_1 _3709_ (.A1(_0908_),
    .A2(_1289_),
    .B1(_0905_),
    .Y(_1290_));
 sky130_fd_sc_hd__o221a_1 _3710_ (.A1(_0905_),
    .A2(_1286_),
    .B1(_1288_),
    .B2(_1290_),
    .C1(net18),
    .X(_1291_));
 sky130_fd_sc_hd__mux4_1 _3711_ (.A0(\dmmu0.page_table[4][12] ),
    .A1(\dmmu0.page_table[5][12] ),
    .A2(\dmmu0.page_table[6][12] ),
    .A3(\dmmu0.page_table[7][12] ),
    .S0(_0895_),
    .S1(net16),
    .X(_1292_));
 sky130_fd_sc_hd__mux2_1 _3712_ (.A0(\dmmu0.page_table[2][12] ),
    .A1(\dmmu0.page_table[3][12] ),
    .S(net15),
    .X(_1293_));
 sky130_fd_sc_hd__mux2_1 _3713_ (.A0(\dmmu0.page_table[0][12] ),
    .A1(\dmmu0.page_table[1][12] ),
    .S(net15),
    .X(_1294_));
 sky130_fd_sc_hd__or2_1 _3714_ (.A(net16),
    .B(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__o211a_1 _3715_ (.A1(_0908_),
    .A2(_1293_),
    .B1(_1295_),
    .C1(_0917_),
    .X(_1296_));
 sky130_fd_sc_hd__a211o_1 _3716_ (.A1(_0905_),
    .A2(_1292_),
    .B1(_1296_),
    .C1(net18),
    .X(_1297_));
 sky130_fd_sc_hd__and3b_1 _3717_ (.A_N(_1291_),
    .B(_1297_),
    .C(_0929_),
    .X(_1298_));
 sky130_fd_sc_hd__a31o_1 _3718_ (.A1(_0957_),
    .A2(_1283_),
    .A3(_1284_),
    .B1(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__o211ai_1 _3719_ (.A1(_1207_),
    .A2(_1208_),
    .B1(_1257_),
    .C1(_1205_),
    .Y(_1300_));
 sky130_fd_sc_hd__xor2_1 _3720_ (.A(net157),
    .B(\dmmu1.long_off_reg[7] ),
    .X(_1301_));
 sky130_fd_sc_hd__a21oi_1 _3721_ (.A1(_1256_),
    .A2(_1300_),
    .B1(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__a31o_1 _3722_ (.A1(_1256_),
    .A2(_1301_),
    .A3(_1300_),
    .B1(_0879_),
    .X(_1303_));
 sky130_fd_sc_hd__mux2_1 _3723_ (.A0(\dmmu1.page_table[2][12] ),
    .A1(\dmmu1.page_table[3][12] ),
    .S(_0857_),
    .X(_1304_));
 sky130_fd_sc_hd__mux2_1 _3724_ (.A0(\dmmu1.page_table[0][12] ),
    .A1(\dmmu1.page_table[1][12] ),
    .S(_1146_),
    .X(_1305_));
 sky130_fd_sc_hd__o21a_1 _3725_ (.A1(_0859_),
    .A2(_1305_),
    .B1(_0871_),
    .X(_1306_));
 sky130_fd_sc_hd__o21ai_1 _3726_ (.A1(_0869_),
    .A2(_1304_),
    .B1(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__mux4_1 _3727_ (.A0(\dmmu1.page_table[4][12] ),
    .A1(\dmmu1.page_table[5][12] ),
    .A2(\dmmu1.page_table[6][12] ),
    .A3(\dmmu1.page_table[7][12] ),
    .S0(_1146_),
    .S1(net121),
    .X(_1308_));
 sky130_fd_sc_hd__a21oi_1 _3728_ (.A1(_0854_),
    .A2(_1308_),
    .B1(net123),
    .Y(_1309_));
 sky130_fd_sc_hd__mux4_1 _3729_ (.A0(\dmmu1.page_table[8][12] ),
    .A1(\dmmu1.page_table[9][12] ),
    .A2(\dmmu1.page_table[10][12] ),
    .A3(\dmmu1.page_table[11][12] ),
    .S0(_1146_),
    .S1(_0859_),
    .X(_1310_));
 sky130_fd_sc_hd__mux2_1 _3730_ (.A0(\dmmu1.page_table[14][12] ),
    .A1(\dmmu1.page_table[15][12] ),
    .S(_0856_),
    .X(_1311_));
 sky130_fd_sc_hd__mux2_1 _3731_ (.A0(\dmmu1.page_table[12][12] ),
    .A1(\dmmu1.page_table[13][12] ),
    .S(net120),
    .X(_1312_));
 sky130_fd_sc_hd__or2_1 _3732_ (.A(net121),
    .B(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__o211a_1 _3733_ (.A1(_0868_),
    .A2(_1311_),
    .B1(_1313_),
    .C1(_0854_),
    .X(_1314_));
 sky130_fd_sc_hd__a211oi_2 _3734_ (.A1(_0872_),
    .A2(_1310_),
    .B1(_1314_),
    .C1(_0874_),
    .Y(_1315_));
 sky130_fd_sc_hd__a21oi_4 _3735_ (.A1(_1307_),
    .A2(_1309_),
    .B1(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__a2bb2o_2 _3736_ (.A1_N(_1302_),
    .A2_N(_1303_),
    .B1(_1316_),
    .B2(_0880_),
    .X(_1317_));
 sky130_fd_sc_hd__mux2_1 _3737_ (.A0(_1299_),
    .A1(_1317_),
    .S(_0818_),
    .X(_1318_));
 sky130_fd_sc_hd__clkbuf_4 _3738_ (.A(_1318_),
    .X(net536));
 sky130_fd_sc_hd__mux2_1 _3739_ (.A0(net134),
    .A1(net29),
    .S(_0847_),
    .X(_1319_));
 sky130_fd_sc_hd__clkbuf_1 _3740_ (.A(_1319_),
    .X(net546));
 sky130_fd_sc_hd__mux2_1 _3741_ (.A0(net141),
    .A1(net36),
    .S(_0847_),
    .X(_1320_));
 sky130_fd_sc_hd__clkbuf_1 _3742_ (.A(_1320_),
    .X(net553));
 sky130_fd_sc_hd__mux2_2 _3743_ (.A0(net142),
    .A1(net37),
    .S(_0847_),
    .X(_1321_));
 sky130_fd_sc_hd__clkbuf_1 _3744_ (.A(_1321_),
    .X(net554));
 sky130_fd_sc_hd__buf_4 _3745_ (.A(_0839_),
    .X(_1322_));
 sky130_fd_sc_hd__mux2_1 _3746_ (.A0(net143),
    .A1(net38),
    .S(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3747_ (.A(_1323_),
    .X(net555));
 sky130_fd_sc_hd__mux2_2 _3748_ (.A0(net144),
    .A1(net39),
    .S(_1322_),
    .X(_1324_));
 sky130_fd_sc_hd__clkbuf_1 _3749_ (.A(_1324_),
    .X(net556));
 sky130_fd_sc_hd__mux2_2 _3750_ (.A0(net145),
    .A1(net40),
    .S(_1322_),
    .X(_1325_));
 sky130_fd_sc_hd__clkbuf_1 _3751_ (.A(_1325_),
    .X(net557));
 sky130_fd_sc_hd__mux2_2 _3752_ (.A0(net146),
    .A1(net41),
    .S(_1322_),
    .X(_1326_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3753_ (.A(_1326_),
    .X(net558));
 sky130_fd_sc_hd__mux2_2 _3754_ (.A0(net147),
    .A1(net42),
    .S(_1322_),
    .X(_1327_));
 sky130_fd_sc_hd__clkbuf_2 _3755_ (.A(_1327_),
    .X(net559));
 sky130_fd_sc_hd__mux2_2 _3756_ (.A0(net148),
    .A1(net43),
    .S(_1322_),
    .X(_1328_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3757_ (.A(_1328_),
    .X(net560));
 sky130_fd_sc_hd__mux2_2 _3758_ (.A0(net149),
    .A1(net44),
    .S(_1322_),
    .X(_1329_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3759_ (.A(_1329_),
    .X(net561));
 sky130_fd_sc_hd__mux2_2 _3760_ (.A0(net135),
    .A1(net30),
    .S(_1322_),
    .X(_1330_));
 sky130_fd_sc_hd__clkbuf_2 _3761_ (.A(_1330_),
    .X(net547));
 sky130_fd_sc_hd__mux2_2 _3762_ (.A0(net136),
    .A1(net31),
    .S(_1322_),
    .X(_1331_));
 sky130_fd_sc_hd__clkbuf_2 _3763_ (.A(_1331_),
    .X(net548));
 sky130_fd_sc_hd__mux2_4 _3764_ (.A0(net137),
    .A1(net32),
    .S(_1322_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_1 _3765_ (.A(_1332_),
    .X(net549));
 sky130_fd_sc_hd__mux2_4 _3766_ (.A0(net138),
    .A1(net33),
    .S(_0839_),
    .X(_1333_));
 sky130_fd_sc_hd__clkbuf_1 _3767_ (.A(_1333_),
    .X(net550));
 sky130_fd_sc_hd__mux2_8 _3768_ (.A0(net139),
    .A1(net34),
    .S(_0839_),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_1 _3769_ (.A(_1334_),
    .X(net551));
 sky130_fd_sc_hd__mux2_8 _3770_ (.A0(net140),
    .A1(net35),
    .S(_0839_),
    .X(_1335_));
 sky130_fd_sc_hd__clkbuf_1 _3771_ (.A(_1335_),
    .X(net552));
 sky130_fd_sc_hd__mux2_1 _3772_ (.A0(net160),
    .A1(net55),
    .S(_0839_),
    .X(_1336_));
 sky130_fd_sc_hd__clkbuf_1 _3773_ (.A(_1336_),
    .X(net563));
 sky130_fd_sc_hd__mux2_1 _3774_ (.A0(net161),
    .A1(net56),
    .S(_0839_),
    .X(_1337_));
 sky130_fd_sc_hd__clkbuf_1 _3775_ (.A(_1337_),
    .X(net564));
 sky130_fd_sc_hd__or3_1 _3776_ (.A(_1194_),
    .B(_1228_),
    .C(_1254_),
    .X(_1338_));
 sky130_fd_sc_hd__or4_1 _3777_ (.A(_0838_),
    .B(_1168_),
    .C(_1211_),
    .D(_1279_),
    .X(_1339_));
 sky130_fd_sc_hd__and3b_2 _3778_ (.A_N(net536),
    .B(_1338_),
    .C(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__clkbuf_1 _3779_ (.A(_1340_),
    .X(net545));
 sky130_fd_sc_hd__and2_1 _3780_ (.A(net212),
    .B(_0993_),
    .X(_1341_));
 sky130_fd_sc_hd__clkbuf_1 _3781_ (.A(_1341_),
    .X(net411));
 sky130_fd_sc_hd__and2_1 _3782_ (.A(net214),
    .B(_0993_),
    .X(_1342_));
 sky130_fd_sc_hd__clkbuf_1 _3783_ (.A(_1342_),
    .X(net412));
 sky130_fd_sc_hd__and2_1 _3784_ (.A(net221),
    .B(_0993_),
    .X(_1343_));
 sky130_fd_sc_hd__clkbuf_1 _3785_ (.A(_1343_),
    .X(net419));
 sky130_fd_sc_hd__and2_1 _3786_ (.A(net222),
    .B(_0993_),
    .X(_1344_));
 sky130_fd_sc_hd__clkbuf_1 _3787_ (.A(_1344_),
    .X(net420));
 sky130_fd_sc_hd__and2_1 _3788_ (.A(net223),
    .B(_0993_),
    .X(_1345_));
 sky130_fd_sc_hd__clkbuf_1 _3789_ (.A(_1345_),
    .X(net421));
 sky130_fd_sc_hd__and2_1 _3790_ (.A(net224),
    .B(_0993_),
    .X(_1346_));
 sky130_fd_sc_hd__clkbuf_1 _3791_ (.A(_1346_),
    .X(net422));
 sky130_fd_sc_hd__and2_1 _3792_ (.A(net225),
    .B(_0993_),
    .X(_1347_));
 sky130_fd_sc_hd__clkbuf_1 _3793_ (.A(_1347_),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 _3794_ (.A(_0839_),
    .X(_1348_));
 sky130_fd_sc_hd__and2_1 _3795_ (.A(net226),
    .B(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__clkbuf_1 _3796_ (.A(_1349_),
    .X(net424));
 sky130_fd_sc_hd__and2_1 _3797_ (.A(net227),
    .B(_1348_),
    .X(_1350_));
 sky130_fd_sc_hd__clkbuf_1 _3798_ (.A(_1350_),
    .X(net425));
 sky130_fd_sc_hd__and2_1 _3799_ (.A(net228),
    .B(_1348_),
    .X(_1351_));
 sky130_fd_sc_hd__clkbuf_1 _3800_ (.A(_1351_),
    .X(net426));
 sky130_fd_sc_hd__and2_1 _3801_ (.A(net229),
    .B(_1348_),
    .X(_1352_));
 sky130_fd_sc_hd__clkbuf_1 _3802_ (.A(_1352_),
    .X(net427));
 sky130_fd_sc_hd__and2_1 _3803_ (.A(net215),
    .B(_1348_),
    .X(_1353_));
 sky130_fd_sc_hd__clkbuf_1 _3804_ (.A(_1353_),
    .X(net413));
 sky130_fd_sc_hd__and2_1 _3805_ (.A(net216),
    .B(_1348_),
    .X(_1354_));
 sky130_fd_sc_hd__clkbuf_1 _3806_ (.A(_1354_),
    .X(net414));
 sky130_fd_sc_hd__and2_1 _3807_ (.A(net217),
    .B(_1348_),
    .X(_1355_));
 sky130_fd_sc_hd__clkbuf_1 _3808_ (.A(_1355_),
    .X(net415));
 sky130_fd_sc_hd__and2_1 _3809_ (.A(net218),
    .B(_1348_),
    .X(_1356_));
 sky130_fd_sc_hd__clkbuf_1 _3810_ (.A(_1356_),
    .X(net416));
 sky130_fd_sc_hd__and2_1 _3811_ (.A(net219),
    .B(_1348_),
    .X(_1357_));
 sky130_fd_sc_hd__clkbuf_1 _3812_ (.A(_1357_),
    .X(net417));
 sky130_fd_sc_hd__and2_1 _3813_ (.A(net220),
    .B(_1348_),
    .X(_1358_));
 sky130_fd_sc_hd__clkbuf_1 _3814_ (.A(_1358_),
    .X(net418));
 sky130_fd_sc_hd__and2_1 _3815_ (.A(net213),
    .B(_0840_),
    .X(_1359_));
 sky130_fd_sc_hd__clkbuf_1 _3816_ (.A(_1359_),
    .X(net428));
 sky130_fd_sc_hd__buf_4 _3817_ (.A(_0812_),
    .X(_1360_));
 sky130_fd_sc_hd__mux2_2 _3818_ (.A0(net328),
    .A1(net382),
    .S(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__mux2_4 _3819_ (.A0(net274),
    .A1(_1361_),
    .S(net664),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_1 _3820_ (.A(_1362_),
    .X(net708));
 sky130_fd_sc_hd__buf_4 _3821_ (.A(\inner_wb_arbiter.o_sel_sig ),
    .X(_1363_));
 sky130_fd_sc_hd__and2_1 _3822_ (.A(_1363_),
    .B(net256),
    .X(_1364_));
 sky130_fd_sc_hd__clkbuf_1 _3823_ (.A(_1364_),
    .X(net690));
 sky130_fd_sc_hd__and2_1 _3824_ (.A(_1363_),
    .B(net263),
    .X(_1365_));
 sky130_fd_sc_hd__clkbuf_1 _3825_ (.A(_1365_),
    .X(net697));
 sky130_fd_sc_hd__and2_1 _3826_ (.A(_1363_),
    .B(net264),
    .X(_1366_));
 sky130_fd_sc_hd__clkbuf_1 _3827_ (.A(_1366_),
    .X(net698));
 sky130_fd_sc_hd__and2_1 _3828_ (.A(_1363_),
    .B(net265),
    .X(_1367_));
 sky130_fd_sc_hd__clkbuf_1 _3829_ (.A(_1367_),
    .X(net699));
 sky130_fd_sc_hd__and2_1 _3830_ (.A(_1363_),
    .B(net266),
    .X(_1368_));
 sky130_fd_sc_hd__clkbuf_1 _3831_ (.A(_1368_),
    .X(net700));
 sky130_fd_sc_hd__and2_1 _3832_ (.A(_1363_),
    .B(net267),
    .X(_1369_));
 sky130_fd_sc_hd__clkbuf_1 _3833_ (.A(_1369_),
    .X(net701));
 sky130_fd_sc_hd__and2_1 _3834_ (.A(_1363_),
    .B(net268),
    .X(_1370_));
 sky130_fd_sc_hd__clkbuf_1 _3835_ (.A(_1370_),
    .X(net702));
 sky130_fd_sc_hd__and2_1 _3836_ (.A(_1363_),
    .B(net269),
    .X(_1371_));
 sky130_fd_sc_hd__clkbuf_1 _3837_ (.A(_1371_),
    .X(net703));
 sky130_fd_sc_hd__and2_1 _3838_ (.A(_1363_),
    .B(net270),
    .X(_1372_));
 sky130_fd_sc_hd__clkbuf_1 _3839_ (.A(_1372_),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_4 _3840_ (.A(\inner_wb_arbiter.o_sel_sig ),
    .X(_1373_));
 sky130_fd_sc_hd__and2_4 _3841_ (.A(_1373_),
    .B(net271),
    .X(_1374_));
 sky130_fd_sc_hd__clkbuf_1 _3842_ (.A(_1374_),
    .X(net705));
 sky130_fd_sc_hd__and2_4 _3843_ (.A(_1373_),
    .B(net257),
    .X(_1375_));
 sky130_fd_sc_hd__clkbuf_1 _3844_ (.A(_1375_),
    .X(net691));
 sky130_fd_sc_hd__and2_4 _3845_ (.A(_1373_),
    .B(net258),
    .X(_1376_));
 sky130_fd_sc_hd__clkbuf_1 _3846_ (.A(_1376_),
    .X(net692));
 sky130_fd_sc_hd__and2_4 _3847_ (.A(_1373_),
    .B(net259),
    .X(_1377_));
 sky130_fd_sc_hd__clkbuf_1 _3848_ (.A(_1377_),
    .X(net693));
 sky130_fd_sc_hd__and2_4 _3849_ (.A(_1373_),
    .B(net260),
    .X(_1378_));
 sky130_fd_sc_hd__clkbuf_1 _3850_ (.A(_1378_),
    .X(net694));
 sky130_fd_sc_hd__and2_4 _3851_ (.A(_1373_),
    .B(net261),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_1 _3852_ (.A(_1379_),
    .X(net695));
 sky130_fd_sc_hd__and2_4 _3853_ (.A(_1373_),
    .B(net262),
    .X(_1380_));
 sky130_fd_sc_hd__clkbuf_1 _3854_ (.A(_1380_),
    .X(net696));
 sky130_fd_sc_hd__mux2_2 _3855_ (.A0(net309),
    .A1(net363),
    .S(_1360_),
    .X(_1381_));
 sky130_fd_sc_hd__mux2_4 _3856_ (.A0(net231),
    .A1(_1381_),
    .S(net664),
    .X(_1382_));
 sky130_fd_sc_hd__clkbuf_1 _3857_ (.A(_1382_),
    .X(net665));
 sky130_fd_sc_hd__mux2_2 _3858_ (.A0(net316),
    .A1(net370),
    .S(_1360_),
    .X(_1383_));
 sky130_fd_sc_hd__mux2_4 _3859_ (.A0(net242),
    .A1(_1383_),
    .S(net664),
    .X(_1384_));
 sky130_fd_sc_hd__clkbuf_1 _3860_ (.A(_1384_),
    .X(net676));
 sky130_fd_sc_hd__mux2_2 _3861_ (.A0(net317),
    .A1(net371),
    .S(_1360_),
    .X(_1385_));
 sky130_fd_sc_hd__buf_6 _3862_ (.A(_0811_),
    .X(_1386_));
 sky130_fd_sc_hd__mux2_4 _3863_ (.A0(net247),
    .A1(_1385_),
    .S(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__clkbuf_1 _3864_ (.A(_1387_),
    .X(net681));
 sky130_fd_sc_hd__mux2_2 _3865_ (.A0(net318),
    .A1(net372),
    .S(_1360_),
    .X(_1388_));
 sky130_fd_sc_hd__mux2_4 _3866_ (.A0(net248),
    .A1(_1388_),
    .S(_1386_),
    .X(_1389_));
 sky130_fd_sc_hd__clkbuf_1 _3867_ (.A(_1389_),
    .X(net682));
 sky130_fd_sc_hd__buf_4 _3868_ (.A(_0812_),
    .X(_1390_));
 sky130_fd_sc_hd__mux2_2 _3869_ (.A0(net319),
    .A1(net373),
    .S(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__mux2_4 _3870_ (.A0(net249),
    .A1(_1391_),
    .S(_1386_),
    .X(_1392_));
 sky130_fd_sc_hd__clkbuf_1 _3871_ (.A(_1392_),
    .X(net683));
 sky130_fd_sc_hd__mux2_2 _3872_ (.A0(net320),
    .A1(net374),
    .S(_1390_),
    .X(_1393_));
 sky130_fd_sc_hd__mux2_4 _3873_ (.A0(net250),
    .A1(_1393_),
    .S(_1386_),
    .X(_1394_));
 sky130_fd_sc_hd__clkbuf_1 _3874_ (.A(_1394_),
    .X(net684));
 sky130_fd_sc_hd__mux2_1 _3875_ (.A0(net321),
    .A1(net375),
    .S(_1390_),
    .X(_1395_));
 sky130_fd_sc_hd__mux2_4 _3876_ (.A0(net251),
    .A1(_1395_),
    .S(_1386_),
    .X(_1396_));
 sky130_fd_sc_hd__clkbuf_1 _3877_ (.A(_1396_),
    .X(net685));
 sky130_fd_sc_hd__mux2_1 _3878_ (.A0(net322),
    .A1(net376),
    .S(_1390_),
    .X(_1397_));
 sky130_fd_sc_hd__mux2_4 _3879_ (.A0(net252),
    .A1(_1397_),
    .S(_1386_),
    .X(_1398_));
 sky130_fd_sc_hd__clkbuf_1 _3880_ (.A(_1398_),
    .X(net686));
 sky130_fd_sc_hd__mux2_1 _3881_ (.A0(net323),
    .A1(net377),
    .S(_1390_),
    .X(_1399_));
 sky130_fd_sc_hd__mux2_4 _3882_ (.A0(net253),
    .A1(_1399_),
    .S(_1386_),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_1 _3883_ (.A(_1400_),
    .X(net687));
 sky130_fd_sc_hd__mux2_1 _3884_ (.A0(net324),
    .A1(net378),
    .S(_1390_),
    .X(_1401_));
 sky130_fd_sc_hd__mux2_4 _3885_ (.A0(net254),
    .A1(_1401_),
    .S(_1386_),
    .X(_1402_));
 sky130_fd_sc_hd__clkbuf_1 _3886_ (.A(_1402_),
    .X(net688));
 sky130_fd_sc_hd__mux2_1 _3887_ (.A0(net310),
    .A1(net364),
    .S(_1390_),
    .X(_1403_));
 sky130_fd_sc_hd__mux2_4 _3888_ (.A0(net232),
    .A1(_1403_),
    .S(_1386_),
    .X(_1404_));
 sky130_fd_sc_hd__clkbuf_1 _3889_ (.A(_1404_),
    .X(net666));
 sky130_fd_sc_hd__mux2_1 _3890_ (.A0(net311),
    .A1(net365),
    .S(_1390_),
    .X(_1405_));
 sky130_fd_sc_hd__mux2_4 _3891_ (.A0(net233),
    .A1(_1405_),
    .S(_1386_),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_1 _3892_ (.A(_1406_),
    .X(net667));
 sky130_fd_sc_hd__buf_6 _3893_ (.A(net312),
    .X(_1407_));
 sky130_fd_sc_hd__clkbuf_8 _3894_ (.A(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__buf_6 _3895_ (.A(_1408_),
    .X(_1409_));
 sky130_fd_sc_hd__nor3b_4 _3896_ (.A(net385),
    .B(net2),
    .C_N(net3),
    .Y(_1410_));
 sky130_fd_sc_hd__clkbuf_4 _3897_ (.A(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__or2_1 _3898_ (.A(_1409_),
    .B(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__clkbuf_4 _3899_ (.A(net315),
    .X(_1413_));
 sky130_fd_sc_hd__mux4_1 _3900_ (.A0(\immu_0.page_table[4][0] ),
    .A1(\immu_0.page_table[5][0] ),
    .A2(\immu_0.page_table[6][0] ),
    .A3(\immu_0.page_table[7][0] ),
    .S0(_1407_),
    .S1(net313),
    .X(_1414_));
 sky130_fd_sc_hd__mux4_1 _3901_ (.A0(\immu_0.page_table[0][0] ),
    .A1(\immu_0.page_table[1][0] ),
    .A2(\immu_0.page_table[2][0] ),
    .A3(\immu_0.page_table[3][0] ),
    .S0(_1407_),
    .S1(net313),
    .X(_1415_));
 sky130_fd_sc_hd__inv_2 _3902_ (.A(net314),
    .Y(_1416_));
 sky130_fd_sc_hd__mux2_1 _3903_ (.A0(_1414_),
    .A1(_1415_),
    .S(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__inv_2 _3904_ (.A(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__buf_4 _3905_ (.A(net313),
    .X(_1419_));
 sky130_fd_sc_hd__buf_4 _3906_ (.A(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__mux2_1 _3907_ (.A0(\immu_0.page_table[14][0] ),
    .A1(\immu_0.page_table[15][0] ),
    .S(_1408_),
    .X(_1421_));
 sky130_fd_sc_hd__nand2_1 _3908_ (.A(_1420_),
    .B(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__clkinv_2 _3909_ (.A(net313),
    .Y(_1423_));
 sky130_fd_sc_hd__clkbuf_4 _3910_ (.A(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__buf_6 _3911_ (.A(_1407_),
    .X(_1425_));
 sky130_fd_sc_hd__mux2_1 _3912_ (.A0(\immu_0.page_table[12][0] ),
    .A1(\immu_0.page_table[13][0] ),
    .S(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__a21oi_1 _3913_ (.A1(_1424_),
    .A2(_1426_),
    .B1(_1416_),
    .Y(_1427_));
 sky130_fd_sc_hd__mux2_1 _3914_ (.A0(\immu_0.page_table[8][0] ),
    .A1(\immu_0.page_table[9][0] ),
    .S(_1408_),
    .X(_1428_));
 sky130_fd_sc_hd__nand2_1 _3915_ (.A(_1424_),
    .B(_1428_),
    .Y(_1429_));
 sky130_fd_sc_hd__buf_4 _3916_ (.A(_1419_),
    .X(_1430_));
 sky130_fd_sc_hd__mux2_1 _3917_ (.A0(\immu_0.page_table[10][0] ),
    .A1(\immu_0.page_table[11][0] ),
    .S(_1425_),
    .X(_1431_));
 sky130_fd_sc_hd__clkbuf_4 _3918_ (.A(net314),
    .X(_1432_));
 sky130_fd_sc_hd__a21oi_1 _3919_ (.A1(_1430_),
    .A2(_1431_),
    .B1(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__inv_2 _3920_ (.A(net315),
    .Y(_1434_));
 sky130_fd_sc_hd__a221o_1 _3921_ (.A1(_1422_),
    .A2(_1427_),
    .B1(_1429_),
    .B2(_1433_),
    .C1(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__o211ai_2 _3922_ (.A1(_1413_),
    .A2(_1418_),
    .B1(_1435_),
    .C1(_1411_),
    .Y(_1436_));
 sky130_fd_sc_hd__buf_6 _3923_ (.A(net366),
    .X(_1437_));
 sky130_fd_sc_hd__buf_6 _3924_ (.A(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__buf_6 _3925_ (.A(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__clkinv_2 _3926_ (.A(net107),
    .Y(_1440_));
 sky130_fd_sc_hd__and3b_2 _3927_ (.A_N(net385),
    .B(net108),
    .C(_1440_),
    .X(_1441_));
 sky130_fd_sc_hd__buf_4 _3928_ (.A(net367),
    .X(_1442_));
 sky130_fd_sc_hd__buf_6 _3929_ (.A(net366),
    .X(_1443_));
 sky130_fd_sc_hd__mux2_1 _3930_ (.A0(\immu_1.page_table[6][0] ),
    .A1(\immu_1.page_table[7][0] ),
    .S(_1443_),
    .X(_1444_));
 sky130_fd_sc_hd__and2_1 _3931_ (.A(_1442_),
    .B(_1444_),
    .X(_1445_));
 sky130_fd_sc_hd__inv_2 _3932_ (.A(net367),
    .Y(_1446_));
 sky130_fd_sc_hd__clkbuf_4 _3933_ (.A(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__buf_4 _3934_ (.A(net366),
    .X(_1448_));
 sky130_fd_sc_hd__mux2_1 _3935_ (.A0(\immu_1.page_table[4][0] ),
    .A1(\immu_1.page_table[5][0] ),
    .S(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__inv_2 _3936_ (.A(net368),
    .Y(_1450_));
 sky130_fd_sc_hd__clkbuf_4 _3937_ (.A(_1450_),
    .X(_1451_));
 sky130_fd_sc_hd__a21o_1 _3938_ (.A1(_1447_),
    .A2(_1449_),
    .B1(_1451_),
    .X(_1452_));
 sky130_fd_sc_hd__buf_6 _3939_ (.A(_1437_),
    .X(_1453_));
 sky130_fd_sc_hd__buf_4 _3940_ (.A(net367),
    .X(_1454_));
 sky130_fd_sc_hd__mux4_1 _3941_ (.A0(\immu_1.page_table[0][0] ),
    .A1(\immu_1.page_table[1][0] ),
    .A2(\immu_1.page_table[2][0] ),
    .A3(\immu_1.page_table[3][0] ),
    .S0(_1453_),
    .S1(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__clkbuf_4 _3942_ (.A(net368),
    .X(_1456_));
 sky130_fd_sc_hd__clkinv_4 _3943_ (.A(net369),
    .Y(_1457_));
 sky130_fd_sc_hd__o221a_1 _3944_ (.A1(_1445_),
    .A2(_1452_),
    .B1(_1455_),
    .B2(_1456_),
    .C1(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__mux4_1 _3945_ (.A0(\immu_1.page_table[12][0] ),
    .A1(\immu_1.page_table[13][0] ),
    .A2(\immu_1.page_table[14][0] ),
    .A3(\immu_1.page_table[15][0] ),
    .S0(_1437_),
    .S1(net367),
    .X(_1459_));
 sky130_fd_sc_hd__mux4_2 _3946_ (.A0(\immu_1.page_table[8][0] ),
    .A1(\immu_1.page_table[9][0] ),
    .A2(\immu_1.page_table[10][0] ),
    .A3(\immu_1.page_table[11][0] ),
    .S0(_1437_),
    .S1(net367),
    .X(_1460_));
 sky130_fd_sc_hd__mux2_1 _3947_ (.A0(_1459_),
    .A1(_1460_),
    .S(_1450_),
    .X(_1461_));
 sky130_fd_sc_hd__or3b_4 _3948_ (.A(net385),
    .B(net107),
    .C_N(net108),
    .X(_1462_));
 sky130_fd_sc_hd__a21o_1 _3949_ (.A1(net369),
    .A2(_1461_),
    .B1(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__o221a_1 _3950_ (.A1(_1439_),
    .A2(_1441_),
    .B1(_1458_),
    .B2(_1463_),
    .C1(_0812_),
    .X(_1464_));
 sky130_fd_sc_hd__a31o_1 _3951_ (.A1(_0813_),
    .A2(_1412_),
    .A3(_1436_),
    .B1(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__mux2_4 _3952_ (.A0(net234),
    .A1(_1465_),
    .S(_0811_),
    .X(_1466_));
 sky130_fd_sc_hd__clkbuf_1 _3953_ (.A(_1466_),
    .X(net668));
 sky130_fd_sc_hd__nand2_1 _3954_ (.A(net313),
    .B(_1416_),
    .Y(_1467_));
 sky130_fd_sc_hd__mux2_1 _3955_ (.A0(\immu_0.page_table[10][1] ),
    .A1(\immu_0.page_table[11][1] ),
    .S(_1425_),
    .X(_1468_));
 sky130_fd_sc_hd__mux4_1 _3956_ (.A0(\immu_0.page_table[12][1] ),
    .A1(\immu_0.page_table[13][1] ),
    .A2(\immu_0.page_table[14][1] ),
    .A3(\immu_0.page_table[15][1] ),
    .S0(net312),
    .S1(net313),
    .X(_1469_));
 sky130_fd_sc_hd__or2_1 _3957_ (.A(_1416_),
    .B(_1469_),
    .X(_1470_));
 sky130_fd_sc_hd__o211a_1 _3958_ (.A1(_1467_),
    .A2(_1468_),
    .B1(net315),
    .C1(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__buf_6 _3959_ (.A(net312),
    .X(_1472_));
 sky130_fd_sc_hd__mux4_2 _3960_ (.A0(\immu_0.page_table[4][1] ),
    .A1(\immu_0.page_table[5][1] ),
    .A2(\immu_0.page_table[6][1] ),
    .A3(\immu_0.page_table[7][1] ),
    .S0(_1472_),
    .S1(_1419_),
    .X(_1473_));
 sky130_fd_sc_hd__mux2_1 _3961_ (.A0(\immu_0.page_table[2][1] ),
    .A1(\immu_0.page_table[3][1] ),
    .S(_1407_),
    .X(_1474_));
 sky130_fd_sc_hd__or2_1 _3962_ (.A(_1467_),
    .B(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__o211a_1 _3963_ (.A1(_1416_),
    .A2(_1473_),
    .B1(_1475_),
    .C1(_1434_),
    .X(_1476_));
 sky130_fd_sc_hd__or3b_2 _3964_ (.A(_1471_),
    .B(_1476_),
    .C_N(_1410_),
    .X(_1477_));
 sky130_fd_sc_hd__clkbuf_4 _3965_ (.A(_1423_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_4 _3966_ (.A(_1432_),
    .X(_1479_));
 sky130_fd_sc_hd__buf_6 _3967_ (.A(_1472_),
    .X(_1480_));
 sky130_fd_sc_hd__mux4_1 _3968_ (.A0(\immu_0.page_table[0][1] ),
    .A1(\immu_0.page_table[1][1] ),
    .A2(\immu_0.page_table[8][1] ),
    .A3(\immu_0.page_table[9][1] ),
    .S0(_1480_),
    .S1(net315),
    .X(_1481_));
 sky130_fd_sc_hd__o21ai_1 _3969_ (.A1(_1479_),
    .A2(_1481_),
    .B1(_1411_),
    .Y(_1482_));
 sky130_fd_sc_hd__nand2_1 _3970_ (.A(_1478_),
    .B(_1482_),
    .Y(_1483_));
 sky130_fd_sc_hd__mux4_1 _3971_ (.A0(\immu_1.page_table[12][1] ),
    .A1(\immu_1.page_table[13][1] ),
    .A2(\immu_1.page_table[14][1] ),
    .A3(\immu_1.page_table[15][1] ),
    .S0(_1453_),
    .S1(_1454_),
    .X(_1484_));
 sky130_fd_sc_hd__mux2_1 _3972_ (.A0(\immu_1.page_table[10][1] ),
    .A1(\immu_1.page_table[11][1] ),
    .S(_1443_),
    .X(_1485_));
 sky130_fd_sc_hd__or3_1 _3973_ (.A(_1447_),
    .B(net368),
    .C(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__o211a_1 _3974_ (.A1(_1451_),
    .A2(_1484_),
    .B1(_1486_),
    .C1(net369),
    .X(_1487_));
 sky130_fd_sc_hd__mux4_1 _3975_ (.A0(\immu_1.page_table[4][1] ),
    .A1(\immu_1.page_table[5][1] ),
    .A2(\immu_1.page_table[6][1] ),
    .A3(\immu_1.page_table[7][1] ),
    .S0(_1437_),
    .S1(net367),
    .X(_1488_));
 sky130_fd_sc_hd__or2_1 _3976_ (.A(_1451_),
    .B(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__mux2_1 _3977_ (.A0(\immu_1.page_table[2][1] ),
    .A1(\immu_1.page_table[3][1] ),
    .S(_1443_),
    .X(_1490_));
 sky130_fd_sc_hd__or3_1 _3978_ (.A(_1447_),
    .B(net368),
    .C(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__a31o_1 _3979_ (.A1(_1457_),
    .A2(_1489_),
    .A3(_1491_),
    .B1(_1462_),
    .X(_1492_));
 sky130_fd_sc_hd__buf_6 _3980_ (.A(_1443_),
    .X(_1493_));
 sky130_fd_sc_hd__mux4_2 _3981_ (.A0(\immu_1.page_table[0][1] ),
    .A1(\immu_1.page_table[1][1] ),
    .A2(\immu_1.page_table[8][1] ),
    .A3(\immu_1.page_table[9][1] ),
    .S0(_1493_),
    .S1(net369),
    .X(_1494_));
 sky130_fd_sc_hd__o21a_1 _3982_ (.A1(_1456_),
    .A2(_1494_),
    .B1(_1441_),
    .X(_1495_));
 sky130_fd_sc_hd__buf_4 _3983_ (.A(_1442_),
    .X(_1496_));
 sky130_fd_sc_hd__o221a_1 _3984_ (.A1(_1487_),
    .A2(_1492_),
    .B1(_1495_),
    .B2(_1496_),
    .C1(_0812_),
    .X(_1497_));
 sky130_fd_sc_hd__a31o_1 _3985_ (.A1(_0813_),
    .A2(_1477_),
    .A3(_1483_),
    .B1(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__mux2_4 _3986_ (.A0(net235),
    .A1(_1498_),
    .S(_0811_),
    .X(_1499_));
 sky130_fd_sc_hd__clkbuf_1 _3987_ (.A(_1499_),
    .X(net669));
 sky130_fd_sc_hd__mux2_1 _3988_ (.A0(\immu_0.page_table[0][2] ),
    .A1(\immu_0.page_table[1][2] ),
    .S(_1480_),
    .X(_1500_));
 sky130_fd_sc_hd__mux2_1 _3989_ (.A0(\immu_0.page_table[2][2] ),
    .A1(\immu_0.page_table[3][2] ),
    .S(_1472_),
    .X(_1501_));
 sky130_fd_sc_hd__a21o_1 _3990_ (.A1(_1419_),
    .A2(_1501_),
    .B1(net315),
    .X(_1502_));
 sky130_fd_sc_hd__a21o_1 _3991_ (.A1(_1478_),
    .A2(_1500_),
    .B1(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__mux2_1 _3992_ (.A0(\immu_0.page_table[10][2] ),
    .A1(\immu_0.page_table[11][2] ),
    .S(_1480_),
    .X(_1504_));
 sky130_fd_sc_hd__mux2_2 _3993_ (.A0(\immu_0.page_table[8][2] ),
    .A1(\immu_0.page_table[9][2] ),
    .S(_1472_),
    .X(_1505_));
 sky130_fd_sc_hd__a21o_1 _3994_ (.A1(_1424_),
    .A2(_1505_),
    .B1(_1434_),
    .X(_1506_));
 sky130_fd_sc_hd__a21o_1 _3995_ (.A1(_1420_),
    .A2(_1504_),
    .B1(_1506_),
    .X(_1507_));
 sky130_fd_sc_hd__a31o_1 _3996_ (.A1(_1411_),
    .A2(_1503_),
    .A3(_1507_),
    .B1(_1479_),
    .X(_1508_));
 sky130_fd_sc_hd__mux4_2 _3997_ (.A0(\immu_0.page_table[4][2] ),
    .A1(\immu_0.page_table[5][2] ),
    .A2(\immu_0.page_table[6][2] ),
    .A3(\immu_0.page_table[7][2] ),
    .S0(_1480_),
    .S1(_1430_),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_1 _3998_ (.A0(\immu_0.page_table[14][2] ),
    .A1(\immu_0.page_table[15][2] ),
    .S(_1408_),
    .X(_1510_));
 sky130_fd_sc_hd__mux2_1 _3999_ (.A0(\immu_0.page_table[12][2] ),
    .A1(\immu_0.page_table[13][2] ),
    .S(_1472_),
    .X(_1511_));
 sky130_fd_sc_hd__or2_1 _4000_ (.A(_1419_),
    .B(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__o211a_1 _4001_ (.A1(_1424_),
    .A2(_1510_),
    .B1(_1512_),
    .C1(net315),
    .X(_1513_));
 sky130_fd_sc_hd__nand2_1 _4002_ (.A(_1432_),
    .B(_1410_),
    .Y(_1514_));
 sky130_fd_sc_hd__a211o_1 _4003_ (.A1(_1434_),
    .A2(_1509_),
    .B1(_1513_),
    .C1(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__clkbuf_4 _4004_ (.A(_1456_),
    .X(_1516_));
 sky130_fd_sc_hd__mux4_1 _4005_ (.A0(\immu_1.page_table[0][2] ),
    .A1(\immu_1.page_table[1][2] ),
    .A2(\immu_1.page_table[2][2] ),
    .A3(\immu_1.page_table[3][2] ),
    .S0(_1453_),
    .S1(_1454_),
    .X(_1517_));
 sky130_fd_sc_hd__or2b_1 _4006_ (.A(\immu_1.page_table[11][2] ),
    .B_N(_1448_),
    .X(_1518_));
 sky130_fd_sc_hd__o21a_1 _4007_ (.A1(_1448_),
    .A2(\immu_1.page_table[10][2] ),
    .B1(_1454_),
    .X(_1519_));
 sky130_fd_sc_hd__mux2_1 _4008_ (.A0(\immu_1.page_table[8][2] ),
    .A1(\immu_1.page_table[9][2] ),
    .S(_1443_),
    .X(_1520_));
 sky130_fd_sc_hd__a221o_2 _4009_ (.A1(_1518_),
    .A2(_1519_),
    .B1(_1520_),
    .B2(_1447_),
    .C1(_1457_),
    .X(_1521_));
 sky130_fd_sc_hd__o211a_1 _4010_ (.A1(net369),
    .A2(_1517_),
    .B1(_1521_),
    .C1(_1441_),
    .X(_1522_));
 sky130_fd_sc_hd__buf_4 _4011_ (.A(_1447_),
    .X(_1523_));
 sky130_fd_sc_hd__buf_6 _4012_ (.A(_1448_),
    .X(_1524_));
 sky130_fd_sc_hd__mux2_1 _4013_ (.A0(\immu_1.page_table[14][2] ),
    .A1(\immu_1.page_table[15][2] ),
    .S(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__mux2_1 _4014_ (.A0(\immu_1.page_table[12][2] ),
    .A1(\immu_1.page_table[13][2] ),
    .S(_1448_),
    .X(_1526_));
 sky130_fd_sc_hd__or2_1 _4015_ (.A(_1442_),
    .B(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__o211a_1 _4016_ (.A1(_1523_),
    .A2(_1525_),
    .B1(_1527_),
    .C1(net369),
    .X(_1528_));
 sky130_fd_sc_hd__mux4_1 _4017_ (.A0(\immu_1.page_table[4][2] ),
    .A1(\immu_1.page_table[5][2] ),
    .A2(\immu_1.page_table[6][2] ),
    .A3(\immu_1.page_table[7][2] ),
    .S0(_1438_),
    .S1(_1442_),
    .X(_1529_));
 sky130_fd_sc_hd__buf_4 _4018_ (.A(_1451_),
    .X(_1530_));
 sky130_fd_sc_hd__a211o_1 _4019_ (.A1(_1457_),
    .A2(_1529_),
    .B1(_1462_),
    .C1(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__o221a_1 _4020_ (.A1(_1516_),
    .A2(_1522_),
    .B1(_1528_),
    .B2(_1531_),
    .C1(_0812_),
    .X(_1532_));
 sky130_fd_sc_hd__a31o_1 _4021_ (.A1(_0813_),
    .A2(_1508_),
    .A3(_1515_),
    .B1(_1532_),
    .X(_1533_));
 sky130_fd_sc_hd__mux2_4 _4022_ (.A0(net236),
    .A1(_1533_),
    .S(_0811_),
    .X(_1534_));
 sky130_fd_sc_hd__clkbuf_1 _4023_ (.A(_1534_),
    .X(net670));
 sky130_fd_sc_hd__buf_2 _4024_ (.A(_1416_),
    .X(_1535_));
 sky130_fd_sc_hd__mux4_1 _4025_ (.A0(\immu_0.page_table[8][3] ),
    .A1(\immu_0.page_table[9][3] ),
    .A2(\immu_0.page_table[10][3] ),
    .A3(\immu_0.page_table[11][3] ),
    .S0(_1472_),
    .S1(_1419_),
    .X(_1536_));
 sky130_fd_sc_hd__and2_1 _4026_ (.A(_1535_),
    .B(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__mux2_1 _4027_ (.A0(\immu_0.page_table[14][3] ),
    .A1(\immu_0.page_table[15][3] ),
    .S(_1408_),
    .X(_1538_));
 sky130_fd_sc_hd__mux2_1 _4028_ (.A0(\immu_0.page_table[12][3] ),
    .A1(\immu_0.page_table[13][3] ),
    .S(_1407_),
    .X(_1539_));
 sky130_fd_sc_hd__or2_1 _4029_ (.A(_1419_),
    .B(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__o211a_1 _4030_ (.A1(_1424_),
    .A2(_1538_),
    .B1(_1540_),
    .C1(_1432_),
    .X(_1541_));
 sky130_fd_sc_hd__nand2_1 _4031_ (.A(_1413_),
    .B(_1410_),
    .Y(_1542_));
 sky130_fd_sc_hd__mux2_1 _4032_ (.A0(\immu_0.page_table[2][3] ),
    .A1(\immu_0.page_table[3][3] ),
    .S(_1472_),
    .X(_1543_));
 sky130_fd_sc_hd__mux2_1 _4033_ (.A0(\immu_0.page_table[0][3] ),
    .A1(\immu_0.page_table[1][3] ),
    .S(net312),
    .X(_1544_));
 sky130_fd_sc_hd__a21o_1 _4034_ (.A1(_1423_),
    .A2(_1544_),
    .B1(_1432_),
    .X(_1545_));
 sky130_fd_sc_hd__a21o_1 _4035_ (.A1(_1419_),
    .A2(_1543_),
    .B1(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__mux2_2 _4036_ (.A0(\immu_0.page_table[4][3] ),
    .A1(\immu_0.page_table[5][3] ),
    .S(_1472_),
    .X(_1547_));
 sky130_fd_sc_hd__mux2_1 _4037_ (.A0(\immu_0.page_table[6][3] ),
    .A1(\immu_0.page_table[7][3] ),
    .S(net312),
    .X(_1548_));
 sky130_fd_sc_hd__a21o_1 _4038_ (.A1(_1419_),
    .A2(_1548_),
    .B1(_1416_),
    .X(_1549_));
 sky130_fd_sc_hd__a21o_1 _4039_ (.A1(_1423_),
    .A2(_1547_),
    .B1(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__a31o_1 _4040_ (.A1(_1410_),
    .A2(_1546_),
    .A3(_1550_),
    .B1(net315),
    .X(_1551_));
 sky130_fd_sc_hd__o31a_2 _4041_ (.A1(_1537_),
    .A2(_1541_),
    .A3(_1542_),
    .B1(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__buf_4 _4042_ (.A(net369),
    .X(_1553_));
 sky130_fd_sc_hd__mux4_1 _4043_ (.A0(\immu_1.page_table[0][3] ),
    .A1(\immu_1.page_table[1][3] ),
    .A2(\immu_1.page_table[2][3] ),
    .A3(\immu_1.page_table[3][3] ),
    .S0(_1453_),
    .S1(_1454_),
    .X(_1554_));
 sky130_fd_sc_hd__or2b_1 _4044_ (.A(\immu_1.page_table[7][3] ),
    .B_N(_1448_),
    .X(_1555_));
 sky130_fd_sc_hd__o21a_1 _4045_ (.A1(_1448_),
    .A2(\immu_1.page_table[6][3] ),
    .B1(net367),
    .X(_1556_));
 sky130_fd_sc_hd__mux2_1 _4046_ (.A0(\immu_1.page_table[4][3] ),
    .A1(\immu_1.page_table[5][3] ),
    .S(_1443_),
    .X(_1557_));
 sky130_fd_sc_hd__a221o_1 _4047_ (.A1(_1555_),
    .A2(_1556_),
    .B1(_1557_),
    .B2(_1447_),
    .C1(_1451_),
    .X(_1558_));
 sky130_fd_sc_hd__o211a_1 _4048_ (.A1(_1456_),
    .A2(_1554_),
    .B1(_1558_),
    .C1(_1441_),
    .X(_1559_));
 sky130_fd_sc_hd__mux2_1 _4049_ (.A0(\immu_1.page_table[14][3] ),
    .A1(\immu_1.page_table[15][3] ),
    .S(_1493_),
    .X(_1560_));
 sky130_fd_sc_hd__mux2_1 _4050_ (.A0(\immu_1.page_table[12][3] ),
    .A1(\immu_1.page_table[13][3] ),
    .S(_1448_),
    .X(_1561_));
 sky130_fd_sc_hd__or2_1 _4051_ (.A(_1442_),
    .B(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__o211a_1 _4052_ (.A1(_1523_),
    .A2(_1560_),
    .B1(_1562_),
    .C1(_1456_),
    .X(_1563_));
 sky130_fd_sc_hd__mux4_2 _4053_ (.A0(\immu_1.page_table[8][3] ),
    .A1(\immu_1.page_table[9][3] ),
    .A2(\immu_1.page_table[10][3] ),
    .A3(\immu_1.page_table[11][3] ),
    .S0(_1438_),
    .S1(_1454_),
    .X(_1564_));
 sky130_fd_sc_hd__a211o_1 _4054_ (.A1(_1530_),
    .A2(_1564_),
    .B1(_1462_),
    .C1(_1457_),
    .X(_1565_));
 sky130_fd_sc_hd__o22a_1 _4055_ (.A1(_1553_),
    .A2(_1559_),
    .B1(_1563_),
    .B2(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__mux2_1 _4056_ (.A0(_1552_),
    .A1(_1566_),
    .S(_1390_),
    .X(_1567_));
 sky130_fd_sc_hd__mux2_1 _4057_ (.A0(net237),
    .A1(_1567_),
    .S(_0811_),
    .X(_1568_));
 sky130_fd_sc_hd__clkbuf_4 _4058_ (.A(_1568_),
    .X(net671));
 sky130_fd_sc_hd__buf_4 _4059_ (.A(\inner_wb_arbiter.o_sel_sig ),
    .X(_1569_));
 sky130_fd_sc_hd__buf_4 _4060_ (.A(_1430_),
    .X(_1570_));
 sky130_fd_sc_hd__mux4_1 _4061_ (.A0(\immu_0.page_table[0][4] ),
    .A1(\immu_0.page_table[1][4] ),
    .A2(\immu_0.page_table[2][4] ),
    .A3(\immu_0.page_table[3][4] ),
    .S0(_1409_),
    .S1(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__mux4_1 _4062_ (.A0(\immu_0.page_table[4][4] ),
    .A1(\immu_0.page_table[5][4] ),
    .A2(\immu_0.page_table[6][4] ),
    .A3(\immu_0.page_table[7][4] ),
    .S0(_1409_),
    .S1(_1420_),
    .X(_1572_));
 sky130_fd_sc_hd__mux4_1 _4063_ (.A0(\immu_0.page_table[8][4] ),
    .A1(\immu_0.page_table[9][4] ),
    .A2(\immu_0.page_table[10][4] ),
    .A3(\immu_0.page_table[11][4] ),
    .S0(_1409_),
    .S1(_1420_),
    .X(_1573_));
 sky130_fd_sc_hd__mux4_1 _4064_ (.A0(\immu_0.page_table[12][4] ),
    .A1(\immu_0.page_table[13][4] ),
    .A2(\immu_0.page_table[14][4] ),
    .A3(\immu_0.page_table[15][4] ),
    .S0(_1409_),
    .S1(_1420_),
    .X(_1574_));
 sky130_fd_sc_hd__mux4_2 _4065_ (.A0(_1571_),
    .A1(_1572_),
    .A2(_1573_),
    .A3(_1574_),
    .S0(_1479_),
    .S1(_1413_),
    .X(_1575_));
 sky130_fd_sc_hd__and2_1 _4066_ (.A(net5),
    .B(\immu_0.high_addr_off[0] ),
    .X(_1576_));
 sky130_fd_sc_hd__o21ai_1 _4067_ (.A1(net5),
    .A2(\immu_0.high_addr_off[0] ),
    .B1(net2),
    .Y(_1577_));
 sky130_fd_sc_hd__nor2_1 _4068_ (.A(_1576_),
    .B(_1577_),
    .Y(_1578_));
 sky130_fd_sc_hd__buf_4 _4069_ (.A(_0812_),
    .X(_1579_));
 sky130_fd_sc_hd__a211o_1 _4070_ (.A1(_1411_),
    .A2(_1575_),
    .B1(_1578_),
    .C1(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__buf_4 _4071_ (.A(_1454_),
    .X(_1581_));
 sky130_fd_sc_hd__mux4_2 _4072_ (.A0(\immu_1.page_table[8][4] ),
    .A1(\immu_1.page_table[9][4] ),
    .A2(\immu_1.page_table[10][4] ),
    .A3(\immu_1.page_table[11][4] ),
    .S0(_1439_),
    .S1(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__mux2_1 _4073_ (.A0(\immu_1.page_table[12][4] ),
    .A1(\immu_1.page_table[13][4] ),
    .S(_1439_),
    .X(_1583_));
 sky130_fd_sc_hd__buf_2 _4074_ (.A(_1446_),
    .X(_1584_));
 sky130_fd_sc_hd__mux2_1 _4075_ (.A0(\immu_1.page_table[14][4] ),
    .A1(\immu_1.page_table[15][4] ),
    .S(_1438_),
    .X(_1585_));
 sky130_fd_sc_hd__or2_1 _4076_ (.A(_1584_),
    .B(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__o211a_1 _4077_ (.A1(_1496_),
    .A2(_1583_),
    .B1(_1586_),
    .C1(_1516_),
    .X(_1587_));
 sky130_fd_sc_hd__a211oi_4 _4078_ (.A1(_1530_),
    .A2(_1582_),
    .B1(_1587_),
    .C1(_1457_),
    .Y(_1588_));
 sky130_fd_sc_hd__mux2_1 _4079_ (.A0(\immu_1.page_table[4][4] ),
    .A1(\immu_1.page_table[5][4] ),
    .S(_1524_),
    .X(_1589_));
 sky130_fd_sc_hd__or2_1 _4080_ (.A(_1496_),
    .B(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__mux2_1 _4081_ (.A0(\immu_1.page_table[6][4] ),
    .A1(\immu_1.page_table[7][4] ),
    .S(_1439_),
    .X(_1591_));
 sky130_fd_sc_hd__o21a_1 _4082_ (.A1(_1523_),
    .A2(_1591_),
    .B1(_1516_),
    .X(_1592_));
 sky130_fd_sc_hd__mux4_1 _4083_ (.A0(\immu_1.page_table[0][4] ),
    .A1(\immu_1.page_table[1][4] ),
    .A2(\immu_1.page_table[2][4] ),
    .A3(\immu_1.page_table[3][4] ),
    .S0(_1439_),
    .S1(_1496_),
    .X(_1593_));
 sky130_fd_sc_hd__a221oi_2 _4084_ (.A1(_1590_),
    .A2(_1592_),
    .B1(_1593_),
    .B2(_1530_),
    .C1(_1553_),
    .Y(_1594_));
 sky130_fd_sc_hd__nor2_1 _4085_ (.A(net110),
    .B(\immu_1.high_addr_off[0] ),
    .Y(_1595_));
 sky130_fd_sc_hd__nand2_1 _4086_ (.A(net110),
    .B(\immu_1.high_addr_off[0] ),
    .Y(_1596_));
 sky130_fd_sc_hd__or3b_1 _4087_ (.A(_1440_),
    .B(_1595_),
    .C_N(_1596_),
    .X(_1597_));
 sky130_fd_sc_hd__o311a_1 _4088_ (.A1(_1462_),
    .A2(_1588_),
    .A3(_1594_),
    .B1(_1597_),
    .C1(_1579_),
    .X(_1598_));
 sky130_fd_sc_hd__nor2_1 _4089_ (.A(_1569_),
    .B(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__a22o_4 _4090_ (.A1(_1569_),
    .A2(net238),
    .B1(_1580_),
    .B2(_1599_),
    .X(net672));
 sky130_fd_sc_hd__mux4_2 _4091_ (.A0(\immu_0.page_table[4][5] ),
    .A1(\immu_0.page_table[5][5] ),
    .A2(\immu_0.page_table[6][5] ),
    .A3(\immu_0.page_table[7][5] ),
    .S0(_1409_),
    .S1(_1570_),
    .X(_1600_));
 sky130_fd_sc_hd__buf_6 _4092_ (.A(_1408_),
    .X(_1601_));
 sky130_fd_sc_hd__mux4_1 _4093_ (.A0(\immu_0.page_table[0][5] ),
    .A1(\immu_0.page_table[1][5] ),
    .A2(\immu_0.page_table[2][5] ),
    .A3(\immu_0.page_table[3][5] ),
    .S0(_1601_),
    .S1(_1420_),
    .X(_1602_));
 sky130_fd_sc_hd__a21o_1 _4094_ (.A1(_1535_),
    .A2(_1602_),
    .B1(_1413_),
    .X(_1603_));
 sky130_fd_sc_hd__a21o_1 _4095_ (.A1(_1479_),
    .A2(_1600_),
    .B1(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__mux4_1 _4096_ (.A0(\immu_0.page_table[12][5] ),
    .A1(\immu_0.page_table[13][5] ),
    .A2(\immu_0.page_table[14][5] ),
    .A3(\immu_0.page_table[15][5] ),
    .S0(_1409_),
    .S1(_1570_),
    .X(_1605_));
 sky130_fd_sc_hd__mux4_1 _4097_ (.A0(\immu_0.page_table[8][5] ),
    .A1(\immu_0.page_table[9][5] ),
    .A2(\immu_0.page_table[10][5] ),
    .A3(\immu_0.page_table[11][5] ),
    .S0(_1601_),
    .S1(_1420_),
    .X(_1606_));
 sky130_fd_sc_hd__a21o_1 _4098_ (.A1(_1535_),
    .A2(_1606_),
    .B1(_1434_),
    .X(_1607_));
 sky130_fd_sc_hd__a21o_1 _4099_ (.A1(_1479_),
    .A2(_1605_),
    .B1(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__nand2_1 _4100_ (.A(net6),
    .B(\immu_0.high_addr_off[1] ),
    .Y(_1609_));
 sky130_fd_sc_hd__or2_1 _4101_ (.A(net6),
    .B(\immu_0.high_addr_off[1] ),
    .X(_1610_));
 sky130_fd_sc_hd__nand3_1 _4102_ (.A(_1576_),
    .B(_1609_),
    .C(_1610_),
    .Y(_1611_));
 sky130_fd_sc_hd__a21o_1 _4103_ (.A1(_1609_),
    .A2(_1610_),
    .B1(_1576_),
    .X(_1612_));
 sky130_fd_sc_hd__a31o_2 _4104_ (.A1(net2),
    .A2(_1611_),
    .A3(_1612_),
    .B1(_1360_),
    .X(_1613_));
 sky130_fd_sc_hd__a31o_1 _4105_ (.A1(_1411_),
    .A2(_1604_),
    .A3(_1608_),
    .B1(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__nand2_1 _4106_ (.A(net111),
    .B(\immu_1.high_addr_off[1] ),
    .Y(_1615_));
 sky130_fd_sc_hd__or2_1 _4107_ (.A(net111),
    .B(\immu_1.high_addr_off[1] ),
    .X(_1616_));
 sky130_fd_sc_hd__and3b_1 _4108_ (.A_N(_1596_),
    .B(_1615_),
    .C(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__a21boi_1 _4109_ (.A1(_1615_),
    .A2(_1616_),
    .B1_N(_1596_),
    .Y(_1618_));
 sky130_fd_sc_hd__mux4_2 _4110_ (.A0(\immu_1.page_table[8][5] ),
    .A1(\immu_1.page_table[9][5] ),
    .A2(\immu_1.page_table[10][5] ),
    .A3(\immu_1.page_table[11][5] ),
    .S0(_1437_),
    .S1(net367),
    .X(_1619_));
 sky130_fd_sc_hd__inv_2 _4111_ (.A(_1619_),
    .Y(_1620_));
 sky130_fd_sc_hd__mux2_1 _4112_ (.A0(\immu_1.page_table[12][5] ),
    .A1(\immu_1.page_table[13][5] ),
    .S(_1493_),
    .X(_1621_));
 sky130_fd_sc_hd__nor2_1 _4113_ (.A(_1581_),
    .B(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__mux2_1 _4114_ (.A0(\immu_1.page_table[14][5] ),
    .A1(\immu_1.page_table[15][5] ),
    .S(_1438_),
    .X(_1623_));
 sky130_fd_sc_hd__o21ai_1 _4115_ (.A1(_1584_),
    .A2(_1623_),
    .B1(_1456_),
    .Y(_1624_));
 sky130_fd_sc_hd__o221a_1 _4116_ (.A1(_1456_),
    .A2(_1620_),
    .B1(_1622_),
    .B2(_1624_),
    .C1(_1553_),
    .X(_1625_));
 sky130_fd_sc_hd__mux2_1 _4117_ (.A0(\immu_1.page_table[0][5] ),
    .A1(\immu_1.page_table[1][5] ),
    .S(_1448_),
    .X(_1626_));
 sky130_fd_sc_hd__or2_1 _4118_ (.A(_1442_),
    .B(_1626_),
    .X(_1627_));
 sky130_fd_sc_hd__mux2_1 _4119_ (.A0(\immu_1.page_table[2][5] ),
    .A1(\immu_1.page_table[3][5] ),
    .S(_1448_),
    .X(_1628_));
 sky130_fd_sc_hd__o21a_1 _4120_ (.A1(_1584_),
    .A2(_1628_),
    .B1(_1451_),
    .X(_1629_));
 sky130_fd_sc_hd__mux4_1 _4121_ (.A0(\immu_1.page_table[4][5] ),
    .A1(\immu_1.page_table[5][5] ),
    .A2(\immu_1.page_table[6][5] ),
    .A3(\immu_1.page_table[7][5] ),
    .S0(_1493_),
    .S1(_1442_),
    .X(_1630_));
 sky130_fd_sc_hd__a221o_1 _4122_ (.A1(_1627_),
    .A2(_1629_),
    .B1(_1630_),
    .B2(_1456_),
    .C1(_1553_),
    .X(_1631_));
 sky130_fd_sc_hd__or3b_1 _4123_ (.A(_1462_),
    .B(_1625_),
    .C_N(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__o311a_2 _4124_ (.A1(_1440_),
    .A2(_1617_),
    .A3(_1618_),
    .B1(_1632_),
    .C1(_1360_),
    .X(_1633_));
 sky130_fd_sc_hd__nor2_1 _4125_ (.A(_1569_),
    .B(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__a22o_4 _4126_ (.A1(_1569_),
    .A2(net239),
    .B1(_1614_),
    .B2(_1634_),
    .X(net673));
 sky130_fd_sc_hd__mux2_1 _4127_ (.A0(\immu_0.page_table[8][6] ),
    .A1(\immu_0.page_table[9][6] ),
    .S(_1601_),
    .X(_1635_));
 sky130_fd_sc_hd__or2_2 _4128_ (.A(_1570_),
    .B(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__mux2_1 _4129_ (.A0(\immu_0.page_table[10][6] ),
    .A1(\immu_0.page_table[11][6] ),
    .S(_1601_),
    .X(_1637_));
 sky130_fd_sc_hd__or2_1 _4130_ (.A(_1478_),
    .B(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__mux4_1 _4131_ (.A0(\immu_0.page_table[12][6] ),
    .A1(\immu_0.page_table[13][6] ),
    .A2(\immu_0.page_table[14][6] ),
    .A3(\immu_0.page_table[15][6] ),
    .S0(_1601_),
    .S1(_1430_),
    .X(_1639_));
 sky130_fd_sc_hd__a21o_1 _4132_ (.A1(_1479_),
    .A2(_1639_),
    .B1(_1434_),
    .X(_1640_));
 sky130_fd_sc_hd__a31o_1 _4133_ (.A1(_1535_),
    .A2(_1636_),
    .A3(_1638_),
    .B1(_1640_),
    .X(_1641_));
 sky130_fd_sc_hd__mux4_2 _4134_ (.A0(\immu_0.page_table[4][6] ),
    .A1(\immu_0.page_table[5][6] ),
    .A2(\immu_0.page_table[6][6] ),
    .A3(\immu_0.page_table[7][6] ),
    .S0(_1409_),
    .S1(_1570_),
    .X(_1642_));
 sky130_fd_sc_hd__mux2_1 _4135_ (.A0(\immu_0.page_table[2][6] ),
    .A1(\immu_0.page_table[3][6] ),
    .S(_1601_),
    .X(_1643_));
 sky130_fd_sc_hd__or2_1 _4136_ (.A(_1478_),
    .B(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__mux2_1 _4137_ (.A0(\immu_0.page_table[0][6] ),
    .A1(\immu_0.page_table[1][6] ),
    .S(_1601_),
    .X(_1645_));
 sky130_fd_sc_hd__o21a_1 _4138_ (.A1(_1570_),
    .A2(_1645_),
    .B1(_1535_),
    .X(_1646_));
 sky130_fd_sc_hd__a221o_1 _4139_ (.A1(_1479_),
    .A2(_1642_),
    .B1(_1644_),
    .B2(_1646_),
    .C1(_1413_),
    .X(_1647_));
 sky130_fd_sc_hd__a21boi_2 _4140_ (.A1(_1576_),
    .A2(_1610_),
    .B1_N(_1609_),
    .Y(_1648_));
 sky130_fd_sc_hd__nor2_1 _4141_ (.A(net7),
    .B(\immu_0.high_addr_off[2] ),
    .Y(_1649_));
 sky130_fd_sc_hd__nand2_1 _4142_ (.A(net7),
    .B(\immu_0.high_addr_off[2] ),
    .Y(_1650_));
 sky130_fd_sc_hd__and2b_1 _4143_ (.A_N(_1649_),
    .B(_1650_),
    .X(_1651_));
 sky130_fd_sc_hd__xnor2_1 _4144_ (.A(_1648_),
    .B(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__a21o_1 _4145_ (.A1(net2),
    .A2(_1652_),
    .B1(_1360_),
    .X(_1653_));
 sky130_fd_sc_hd__a31o_1 _4146_ (.A1(_1411_),
    .A2(_1641_),
    .A3(_1647_),
    .B1(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__mux2_1 _4147_ (.A0(\immu_1.page_table[12][6] ),
    .A1(\immu_1.page_table[13][6] ),
    .S(_1453_),
    .X(_1655_));
 sky130_fd_sc_hd__mux2_1 _4148_ (.A0(\immu_1.page_table[14][6] ),
    .A1(\immu_1.page_table[15][6] ),
    .S(_1437_),
    .X(_1656_));
 sky130_fd_sc_hd__or2_1 _4149_ (.A(_1447_),
    .B(_1656_),
    .X(_1657_));
 sky130_fd_sc_hd__o211a_1 _4150_ (.A1(_1442_),
    .A2(_1655_),
    .B1(_1657_),
    .C1(_1456_),
    .X(_1658_));
 sky130_fd_sc_hd__mux2_1 _4151_ (.A0(\immu_1.page_table[10][6] ),
    .A1(\immu_1.page_table[11][6] ),
    .S(_1453_),
    .X(_1659_));
 sky130_fd_sc_hd__mux2_1 _4152_ (.A0(\immu_1.page_table[8][6] ),
    .A1(\immu_1.page_table[9][6] ),
    .S(_1437_),
    .X(_1660_));
 sky130_fd_sc_hd__or2_1 _4153_ (.A(_1454_),
    .B(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__o211a_1 _4154_ (.A1(_1584_),
    .A2(_1659_),
    .B1(_1661_),
    .C1(_1451_),
    .X(_1662_));
 sky130_fd_sc_hd__or3_1 _4155_ (.A(_1457_),
    .B(_1658_),
    .C(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__mux2_1 _4156_ (.A0(\immu_1.page_table[4][6] ),
    .A1(\immu_1.page_table[5][6] ),
    .S(_1438_),
    .X(_1664_));
 sky130_fd_sc_hd__or2_1 _4157_ (.A(_1581_),
    .B(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__mux2_1 _4158_ (.A0(\immu_1.page_table[6][6] ),
    .A1(\immu_1.page_table[7][6] ),
    .S(_1453_),
    .X(_1666_));
 sky130_fd_sc_hd__or2_1 _4159_ (.A(_1584_),
    .B(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__mux2_1 _4160_ (.A0(\immu_1.page_table[0][6] ),
    .A1(\immu_1.page_table[1][6] ),
    .S(_1438_),
    .X(_1668_));
 sky130_fd_sc_hd__mux2_1 _4161_ (.A0(\immu_1.page_table[2][6] ),
    .A1(\immu_1.page_table[3][6] ),
    .S(_1437_),
    .X(_1669_));
 sky130_fd_sc_hd__or2_1 _4162_ (.A(_1447_),
    .B(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__o211a_1 _4163_ (.A1(_1581_),
    .A2(_1668_),
    .B1(_1670_),
    .C1(_1451_),
    .X(_1671_));
 sky130_fd_sc_hd__a311o_1 _4164_ (.A1(_1516_),
    .A2(_1665_),
    .A3(_1667_),
    .B1(_1671_),
    .C1(_1553_),
    .X(_1672_));
 sky130_fd_sc_hd__and3_1 _4165_ (.A(_1441_),
    .B(_1663_),
    .C(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__nor2_1 _4166_ (.A(net111),
    .B(\immu_1.high_addr_off[1] ),
    .Y(_1674_));
 sky130_fd_sc_hd__o21a_1 _4167_ (.A1(_1596_),
    .A2(_1674_),
    .B1(_1615_),
    .X(_1675_));
 sky130_fd_sc_hd__nor2_1 _4168_ (.A(net112),
    .B(\immu_1.high_addr_off[2] ),
    .Y(_1676_));
 sky130_fd_sc_hd__nand2_1 _4169_ (.A(net112),
    .B(\immu_1.high_addr_off[2] ),
    .Y(_1677_));
 sky130_fd_sc_hd__and2b_1 _4170_ (.A_N(_1676_),
    .B(_1677_),
    .X(_1678_));
 sky130_fd_sc_hd__xor2_1 _4171_ (.A(_1675_),
    .B(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__nor2_1 _4172_ (.A(_1440_),
    .B(_1679_),
    .Y(_1680_));
 sky130_fd_sc_hd__o31a_2 _4173_ (.A1(_0813_),
    .A2(_1673_),
    .A3(_1680_),
    .B1(net664),
    .X(_1681_));
 sky130_fd_sc_hd__a22o_4 _4174_ (.A1(_1569_),
    .A2(net240),
    .B1(_1654_),
    .B2(_1681_),
    .X(net674));
 sky130_fd_sc_hd__o211a_1 _4175_ (.A1(_1596_),
    .A2(_1674_),
    .B1(_1677_),
    .C1(_1615_),
    .X(_1682_));
 sky130_fd_sc_hd__nand2_1 _4176_ (.A(net113),
    .B(\immu_1.high_addr_off[3] ),
    .Y(_1683_));
 sky130_fd_sc_hd__or2_1 _4177_ (.A(net113),
    .B(\immu_1.high_addr_off[3] ),
    .X(_1684_));
 sky130_fd_sc_hd__nand2_1 _4178_ (.A(_1683_),
    .B(_1684_),
    .Y(_1685_));
 sky130_fd_sc_hd__o21a_1 _4179_ (.A1(_1676_),
    .A2(_1682_),
    .B1(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__o31ai_1 _4180_ (.A1(_1676_),
    .A2(_1685_),
    .A3(_1682_),
    .B1(net107),
    .Y(_1687_));
 sky130_fd_sc_hd__mux2_1 _4181_ (.A0(\immu_1.page_table[2][7] ),
    .A1(\immu_1.page_table[3][7] ),
    .S(_1493_),
    .X(_1688_));
 sky130_fd_sc_hd__mux2_1 _4182_ (.A0(\immu_1.page_table[0][7] ),
    .A1(\immu_1.page_table[1][7] ),
    .S(_1443_),
    .X(_1689_));
 sky130_fd_sc_hd__or2_1 _4183_ (.A(_1442_),
    .B(_1689_),
    .X(_1690_));
 sky130_fd_sc_hd__o211a_1 _4184_ (.A1(_1523_),
    .A2(_1688_),
    .B1(_1690_),
    .C1(_1530_),
    .X(_1691_));
 sky130_fd_sc_hd__mux2_1 _4185_ (.A0(\immu_1.page_table[4][7] ),
    .A1(\immu_1.page_table[5][7] ),
    .S(_1493_),
    .X(_1692_));
 sky130_fd_sc_hd__mux2_1 _4186_ (.A0(\immu_1.page_table[6][7] ),
    .A1(\immu_1.page_table[7][7] ),
    .S(_1443_),
    .X(_1693_));
 sky130_fd_sc_hd__or2_1 _4187_ (.A(_1447_),
    .B(_1693_),
    .X(_1694_));
 sky130_fd_sc_hd__o211a_1 _4188_ (.A1(_1581_),
    .A2(_1692_),
    .B1(_1694_),
    .C1(_1456_),
    .X(_1695_));
 sky130_fd_sc_hd__mux2_1 _4189_ (.A0(\immu_1.page_table[8][7] ),
    .A1(\immu_1.page_table[9][7] ),
    .S(_1443_),
    .X(_1696_));
 sky130_fd_sc_hd__mux2_1 _4190_ (.A0(\immu_1.page_table[10][7] ),
    .A1(\immu_1.page_table[11][7] ),
    .S(net366),
    .X(_1697_));
 sky130_fd_sc_hd__or2_1 _4191_ (.A(_1446_),
    .B(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__o211a_1 _4192_ (.A1(_1454_),
    .A2(_1696_),
    .B1(_1698_),
    .C1(_1451_),
    .X(_1699_));
 sky130_fd_sc_hd__mux2_1 _4193_ (.A0(\immu_1.page_table[12][7] ),
    .A1(\immu_1.page_table[13][7] ),
    .S(_1443_),
    .X(_1700_));
 sky130_fd_sc_hd__mux2_1 _4194_ (.A0(\immu_1.page_table[14][7] ),
    .A1(\immu_1.page_table[15][7] ),
    .S(net366),
    .X(_1701_));
 sky130_fd_sc_hd__or2_1 _4195_ (.A(_1446_),
    .B(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__o211a_1 _4196_ (.A1(_1454_),
    .A2(_1700_),
    .B1(_1702_),
    .C1(net368),
    .X(_1703_));
 sky130_fd_sc_hd__or3_2 _4197_ (.A(_1457_),
    .B(_1699_),
    .C(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__o31ai_1 _4198_ (.A1(_1553_),
    .A2(_1691_),
    .A3(_1695_),
    .B1(_1704_),
    .Y(_1705_));
 sky130_fd_sc_hd__o221a_1 _4199_ (.A1(_1686_),
    .A2(_1687_),
    .B1(_1705_),
    .B2(_1462_),
    .C1(_1360_),
    .X(_1706_));
 sky130_fd_sc_hd__nand2_1 _4200_ (.A(net8),
    .B(\immu_0.high_addr_off[3] ),
    .Y(_1707_));
 sky130_fd_sc_hd__or2_1 _4201_ (.A(net8),
    .B(\immu_0.high_addr_off[3] ),
    .X(_1708_));
 sky130_fd_sc_hd__o21ai_2 _4202_ (.A1(_1648_),
    .A2(_1649_),
    .B1(_1650_),
    .Y(_1709_));
 sky130_fd_sc_hd__a21o_1 _4203_ (.A1(_1707_),
    .A2(_1708_),
    .B1(_1709_),
    .X(_1710_));
 sky130_fd_sc_hd__nand3_1 _4204_ (.A(_1707_),
    .B(_1708_),
    .C(_1709_),
    .Y(_1711_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(\immu_0.page_table[4][7] ),
    .A1(\immu_0.page_table[5][7] ),
    .S(_1472_),
    .X(_1712_));
 sky130_fd_sc_hd__mux2_1 _4206_ (.A0(\immu_0.page_table[6][7] ),
    .A1(\immu_0.page_table[7][7] ),
    .S(net312),
    .X(_1713_));
 sky130_fd_sc_hd__or2_1 _4207_ (.A(_1423_),
    .B(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__o211a_1 _4208_ (.A1(_1430_),
    .A2(_1712_),
    .B1(_1714_),
    .C1(_1432_),
    .X(_1715_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(\immu_0.page_table[0][7] ),
    .A1(\immu_0.page_table[1][7] ),
    .S(_1425_),
    .X(_1716_));
 sky130_fd_sc_hd__mux2_1 _4210_ (.A0(\immu_0.page_table[2][7] ),
    .A1(\immu_0.page_table[3][7] ),
    .S(net312),
    .X(_1717_));
 sky130_fd_sc_hd__or2_1 _4211_ (.A(_1423_),
    .B(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__o211a_1 _4212_ (.A1(_1430_),
    .A2(_1716_),
    .B1(_1718_),
    .C1(_1416_),
    .X(_1719_));
 sky130_fd_sc_hd__mux2_1 _4213_ (.A0(\immu_0.page_table[14][7] ),
    .A1(\immu_0.page_table[15][7] ),
    .S(_1407_),
    .X(_1720_));
 sky130_fd_sc_hd__mux2_1 _4214_ (.A0(\immu_0.page_table[12][7] ),
    .A1(\immu_0.page_table[13][7] ),
    .S(net312),
    .X(_1721_));
 sky130_fd_sc_hd__or2_1 _4215_ (.A(net313),
    .B(_1721_),
    .X(_1722_));
 sky130_fd_sc_hd__o211a_1 _4216_ (.A1(_1423_),
    .A2(_1720_),
    .B1(_1722_),
    .C1(_1432_),
    .X(_1723_));
 sky130_fd_sc_hd__mux2_1 _4217_ (.A0(\immu_0.page_table[10][7] ),
    .A1(\immu_0.page_table[11][7] ),
    .S(_1407_),
    .X(_1724_));
 sky130_fd_sc_hd__mux2_1 _4218_ (.A0(\immu_0.page_table[8][7] ),
    .A1(\immu_0.page_table[9][7] ),
    .S(net312),
    .X(_1725_));
 sky130_fd_sc_hd__or2_1 _4219_ (.A(net313),
    .B(_1725_),
    .X(_1726_));
 sky130_fd_sc_hd__o211a_1 _4220_ (.A1(_1423_),
    .A2(_1724_),
    .B1(_1726_),
    .C1(_1416_),
    .X(_1727_));
 sky130_fd_sc_hd__o31a_1 _4221_ (.A1(_1434_),
    .A2(_1723_),
    .A3(_1727_),
    .B1(_1410_),
    .X(_1728_));
 sky130_fd_sc_hd__o31a_1 _4222_ (.A1(_1413_),
    .A2(_1715_),
    .A3(_1719_),
    .B1(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__a311o_1 _4223_ (.A1(net2),
    .A2(_1710_),
    .A3(_1711_),
    .B1(_1729_),
    .C1(_0812_),
    .X(_1730_));
 sky130_fd_sc_hd__or3b_1 _4224_ (.A(\inner_wb_arbiter.o_sel_sig ),
    .B(_1706_),
    .C_N(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__a21bo_4 _4225_ (.A1(_1569_),
    .A2(net241),
    .B1_N(_1731_),
    .X(net675));
 sky130_fd_sc_hd__and2_1 _4226_ (.A(net9),
    .B(\immu_0.high_addr_off[4] ),
    .X(_1732_));
 sky130_fd_sc_hd__nor2_1 _4227_ (.A(net9),
    .B(\immu_0.high_addr_off[4] ),
    .Y(_1733_));
 sky130_fd_sc_hd__nor2_1 _4228_ (.A(_1732_),
    .B(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__a21boi_2 _4229_ (.A1(_1708_),
    .A2(_1709_),
    .B1_N(_1707_),
    .Y(_1735_));
 sky130_fd_sc_hd__xnor2_2 _4230_ (.A(_1734_),
    .B(_1735_),
    .Y(_1736_));
 sky130_fd_sc_hd__mux2_1 _4231_ (.A0(\immu_0.page_table[4][8] ),
    .A1(\immu_0.page_table[5][8] ),
    .S(_1601_),
    .X(_1737_));
 sky130_fd_sc_hd__mux2_1 _4232_ (.A0(\immu_0.page_table[6][8] ),
    .A1(\immu_0.page_table[7][8] ),
    .S(_1408_),
    .X(_1738_));
 sky130_fd_sc_hd__or2_1 _4233_ (.A(_1424_),
    .B(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__o211a_1 _4234_ (.A1(_1570_),
    .A2(_1737_),
    .B1(_1739_),
    .C1(_1479_),
    .X(_1740_));
 sky130_fd_sc_hd__mux2_1 _4235_ (.A0(\immu_0.page_table[0][8] ),
    .A1(\immu_0.page_table[1][8] ),
    .S(_1409_),
    .X(_1741_));
 sky130_fd_sc_hd__mux2_1 _4236_ (.A0(\immu_0.page_table[2][8] ),
    .A1(\immu_0.page_table[3][8] ),
    .S(_1408_),
    .X(_1742_));
 sky130_fd_sc_hd__or2_1 _4237_ (.A(_1478_),
    .B(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__o211a_1 _4238_ (.A1(_1570_),
    .A2(_1741_),
    .B1(_1743_),
    .C1(_1535_),
    .X(_1744_));
 sky130_fd_sc_hd__mux2_1 _4239_ (.A0(\immu_0.page_table[10][8] ),
    .A1(\immu_0.page_table[11][8] ),
    .S(_1409_),
    .X(_1745_));
 sky130_fd_sc_hd__mux2_1 _4240_ (.A0(\immu_0.page_table[8][8] ),
    .A1(\immu_0.page_table[9][8] ),
    .S(_1480_),
    .X(_1746_));
 sky130_fd_sc_hd__or2_1 _4241_ (.A(_1420_),
    .B(_1746_),
    .X(_1747_));
 sky130_fd_sc_hd__o211a_1 _4242_ (.A1(_1478_),
    .A2(_1745_),
    .B1(_1747_),
    .C1(_1535_),
    .X(_1748_));
 sky130_fd_sc_hd__mux2_1 _4243_ (.A0(\immu_0.page_table[12][8] ),
    .A1(\immu_0.page_table[13][8] ),
    .S(_1480_),
    .X(_1749_));
 sky130_fd_sc_hd__or2_1 _4244_ (.A(_1420_),
    .B(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__mux2_1 _4245_ (.A0(\immu_0.page_table[14][8] ),
    .A1(\immu_0.page_table[15][8] ),
    .S(_1480_),
    .X(_1751_));
 sky130_fd_sc_hd__or2_1 _4246_ (.A(_1478_),
    .B(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__a31o_1 _4247_ (.A1(_1479_),
    .A2(_1750_),
    .A3(_1752_),
    .B1(_1434_),
    .X(_1753_));
 sky130_fd_sc_hd__o32a_2 _4248_ (.A1(_1413_),
    .A2(_1740_),
    .A3(_1744_),
    .B1(_1748_),
    .B2(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__a221oi_4 _4249_ (.A1(net2),
    .A2(_1736_),
    .B1(_1754_),
    .B2(_1411_),
    .C1(_1579_),
    .Y(_1755_));
 sky130_fd_sc_hd__nand2_1 _4250_ (.A(net114),
    .B(\immu_1.high_addr_off[4] ),
    .Y(_1756_));
 sky130_fd_sc_hd__o21ai_1 _4251_ (.A1(_1676_),
    .A2(_1682_),
    .B1(_1683_),
    .Y(_1757_));
 sky130_fd_sc_hd__or2_1 _4252_ (.A(net114),
    .B(\immu_1.high_addr_off[4] ),
    .X(_1758_));
 sky130_fd_sc_hd__and3_1 _4253_ (.A(_1684_),
    .B(_1757_),
    .C(_1758_),
    .X(_1759_));
 sky130_fd_sc_hd__a22oi_1 _4254_ (.A1(_1684_),
    .A2(_1757_),
    .B1(_1758_),
    .B2(_1756_),
    .Y(_1760_));
 sky130_fd_sc_hd__a211o_1 _4255_ (.A1(_1756_),
    .A2(_1759_),
    .B1(_1760_),
    .C1(_1440_),
    .X(_1761_));
 sky130_fd_sc_hd__mux2_1 _4256_ (.A0(\immu_1.page_table[8][8] ),
    .A1(\immu_1.page_table[9][8] ),
    .S(_1524_),
    .X(_1762_));
 sky130_fd_sc_hd__nor2_1 _4257_ (.A(_1581_),
    .B(_1762_),
    .Y(_1763_));
 sky130_fd_sc_hd__mux2_1 _4258_ (.A0(\immu_1.page_table[10][8] ),
    .A1(\immu_1.page_table[11][8] ),
    .S(_1493_),
    .X(_1764_));
 sky130_fd_sc_hd__o21ai_1 _4259_ (.A1(_1523_),
    .A2(_1764_),
    .B1(_1530_),
    .Y(_1765_));
 sky130_fd_sc_hd__mux2_1 _4260_ (.A0(\immu_1.page_table[14][8] ),
    .A1(\immu_1.page_table[15][8] ),
    .S(_1524_),
    .X(_1766_));
 sky130_fd_sc_hd__nor2_1 _4261_ (.A(_1523_),
    .B(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hd__mux2_1 _4262_ (.A0(\immu_1.page_table[12][8] ),
    .A1(\immu_1.page_table[13][8] ),
    .S(_1524_),
    .X(_1768_));
 sky130_fd_sc_hd__o21ai_1 _4263_ (.A1(_1581_),
    .A2(_1768_),
    .B1(_1516_),
    .Y(_1769_));
 sky130_fd_sc_hd__o221a_2 _4264_ (.A1(_1763_),
    .A2(_1765_),
    .B1(_1767_),
    .B2(_1769_),
    .C1(_1553_),
    .X(_1770_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(\immu_1.page_table[6][8] ),
    .A1(\immu_1.page_table[7][8] ),
    .S(_1453_),
    .X(_1771_));
 sky130_fd_sc_hd__or2_1 _4266_ (.A(_1584_),
    .B(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__mux2_1 _4267_ (.A0(\immu_1.page_table[4][8] ),
    .A1(\immu_1.page_table[5][8] ),
    .S(_1453_),
    .X(_1773_));
 sky130_fd_sc_hd__or2_1 _4268_ (.A(_1442_),
    .B(_1773_),
    .X(_1774_));
 sky130_fd_sc_hd__mux2_1 _4269_ (.A0(\immu_1.page_table[0][8] ),
    .A1(\immu_1.page_table[1][8] ),
    .S(_1438_),
    .X(_1775_));
 sky130_fd_sc_hd__mux2_1 _4270_ (.A0(\immu_1.page_table[2][8] ),
    .A1(\immu_1.page_table[3][8] ),
    .S(_1437_),
    .X(_1776_));
 sky130_fd_sc_hd__or2_1 _4271_ (.A(_1447_),
    .B(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__o211a_1 _4272_ (.A1(_1581_),
    .A2(_1775_),
    .B1(_1777_),
    .C1(_1451_),
    .X(_1778_));
 sky130_fd_sc_hd__a311o_1 _4273_ (.A1(_1516_),
    .A2(_1772_),
    .A3(_1774_),
    .B1(_1778_),
    .C1(_1553_),
    .X(_1779_));
 sky130_fd_sc_hd__or3b_1 _4274_ (.A(_1462_),
    .B(_1770_),
    .C_N(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__a31o_1 _4275_ (.A1(_1579_),
    .A2(_1761_),
    .A3(_1780_),
    .B1(\inner_wb_arbiter.o_sel_sig ),
    .X(_1781_));
 sky130_fd_sc_hd__a2bb2o_4 _4276_ (.A1_N(_1755_),
    .A2_N(_1781_),
    .B1(_1569_),
    .B2(net243),
    .X(net677));
 sky130_fd_sc_hd__and2_1 _4277_ (.A(net10),
    .B(\immu_0.high_addr_off[5] ),
    .X(_1782_));
 sky130_fd_sc_hd__or2_1 _4278_ (.A(net10),
    .B(\immu_0.high_addr_off[5] ),
    .X(_1783_));
 sky130_fd_sc_hd__or2b_1 _4279_ (.A(_1782_),
    .B_N(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__o21bai_1 _4280_ (.A1(_1733_),
    .A2(_1735_),
    .B1_N(_1732_),
    .Y(_1785_));
 sky130_fd_sc_hd__xnor2_1 _4281_ (.A(_1784_),
    .B(_1785_),
    .Y(_1786_));
 sky130_fd_sc_hd__mux2_1 _4282_ (.A0(\immu_0.page_table[6][9] ),
    .A1(\immu_0.page_table[7][9] ),
    .S(_1601_),
    .X(_1787_));
 sky130_fd_sc_hd__mux2_1 _4283_ (.A0(\immu_0.page_table[4][9] ),
    .A1(\immu_0.page_table[5][9] ),
    .S(_1425_),
    .X(_1788_));
 sky130_fd_sc_hd__or2_1 _4284_ (.A(_1430_),
    .B(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__o211a_1 _4285_ (.A1(_1478_),
    .A2(_1787_),
    .B1(_1789_),
    .C1(_1479_),
    .X(_1790_));
 sky130_fd_sc_hd__mux2_1 _4286_ (.A0(\immu_0.page_table[0][9] ),
    .A1(\immu_0.page_table[1][9] ),
    .S(_1601_),
    .X(_1791_));
 sky130_fd_sc_hd__mux2_1 _4287_ (.A0(\immu_0.page_table[2][9] ),
    .A1(\immu_0.page_table[3][9] ),
    .S(_1425_),
    .X(_1792_));
 sky130_fd_sc_hd__or2_1 _4288_ (.A(_1424_),
    .B(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__o211a_1 _4289_ (.A1(_1570_),
    .A2(_1791_),
    .B1(_1793_),
    .C1(_1535_),
    .X(_1794_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(\immu_0.page_table[8][9] ),
    .A1(\immu_0.page_table[9][9] ),
    .S(_1425_),
    .X(_1795_));
 sky130_fd_sc_hd__or2_1 _4291_ (.A(_1430_),
    .B(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__mux2_1 _4292_ (.A0(\immu_0.page_table[10][9] ),
    .A1(\immu_0.page_table[11][9] ),
    .S(_1425_),
    .X(_1797_));
 sky130_fd_sc_hd__or2_1 _4293_ (.A(_1424_),
    .B(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__mux2_1 _4294_ (.A0(\immu_0.page_table[14][9] ),
    .A1(\immu_0.page_table[15][9] ),
    .S(_1408_),
    .X(_1799_));
 sky130_fd_sc_hd__mux2_1 _4295_ (.A0(\immu_0.page_table[12][9] ),
    .A1(\immu_0.page_table[13][9] ),
    .S(_1407_),
    .X(_1800_));
 sky130_fd_sc_hd__or2_1 _4296_ (.A(_1419_),
    .B(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__o211a_1 _4297_ (.A1(_1424_),
    .A2(_1799_),
    .B1(_1801_),
    .C1(_1432_),
    .X(_1802_));
 sky130_fd_sc_hd__a311o_1 _4298_ (.A1(_1535_),
    .A2(_1796_),
    .A3(_1798_),
    .B1(_1434_),
    .C1(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__o31a_1 _4299_ (.A1(_1413_),
    .A2(_1790_),
    .A3(_1794_),
    .B1(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__a221o_1 _4300_ (.A1(net2),
    .A2(_1786_),
    .B1(_1804_),
    .B2(_1411_),
    .C1(_1579_),
    .X(_1805_));
 sky130_fd_sc_hd__and2_1 _4301_ (.A(net115),
    .B(\immu_1.high_addr_off[5] ),
    .X(_1806_));
 sky130_fd_sc_hd__or2_1 _4302_ (.A(net115),
    .B(\immu_1.high_addr_off[5] ),
    .X(_1807_));
 sky130_fd_sc_hd__or2b_1 _4303_ (.A(_1806_),
    .B_N(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__a21o_1 _4304_ (.A1(net114),
    .A2(\immu_1.high_addr_off[4] ),
    .B1(_1759_),
    .X(_1809_));
 sky130_fd_sc_hd__xnor2_1 _4305_ (.A(_1808_),
    .B(_1809_),
    .Y(_1810_));
 sky130_fd_sc_hd__mux2_1 _4306_ (.A0(\immu_1.page_table[12][9] ),
    .A1(\immu_1.page_table[13][9] ),
    .S(_1524_),
    .X(_1811_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(\immu_1.page_table[14][9] ),
    .A1(\immu_1.page_table[15][9] ),
    .S(_1453_),
    .X(_1812_));
 sky130_fd_sc_hd__or2_1 _4308_ (.A(_1584_),
    .B(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__o211a_1 _4309_ (.A1(_1496_),
    .A2(_1811_),
    .B1(_1813_),
    .C1(_1516_),
    .X(_1814_));
 sky130_fd_sc_hd__mux2_1 _4310_ (.A0(\immu_1.page_table[10][9] ),
    .A1(\immu_1.page_table[11][9] ),
    .S(_1524_),
    .X(_1815_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(\immu_1.page_table[8][9] ),
    .A1(\immu_1.page_table[9][9] ),
    .S(_1438_),
    .X(_1816_));
 sky130_fd_sc_hd__or2_1 _4312_ (.A(_1581_),
    .B(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__o211a_1 _4313_ (.A1(_1523_),
    .A2(_1815_),
    .B1(_1817_),
    .C1(_1530_),
    .X(_1818_));
 sky130_fd_sc_hd__mux2_1 _4314_ (.A0(\immu_1.page_table[4][9] ),
    .A1(\immu_1.page_table[5][9] ),
    .S(_1439_),
    .X(_1819_));
 sky130_fd_sc_hd__mux2_1 _4315_ (.A0(\immu_1.page_table[6][9] ),
    .A1(\immu_1.page_table[7][9] ),
    .S(_1493_),
    .X(_1820_));
 sky130_fd_sc_hd__or2_1 _4316_ (.A(_1584_),
    .B(_1820_),
    .X(_1821_));
 sky130_fd_sc_hd__o211a_1 _4317_ (.A1(_1496_),
    .A2(_1819_),
    .B1(_1821_),
    .C1(_1516_),
    .X(_1822_));
 sky130_fd_sc_hd__mux2_1 _4318_ (.A0(\immu_1.page_table[2][9] ),
    .A1(\immu_1.page_table[3][9] ),
    .S(_1493_),
    .X(_1823_));
 sky130_fd_sc_hd__or2_1 _4319_ (.A(_1584_),
    .B(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__mux2_1 _4320_ (.A0(\immu_1.page_table[0][9] ),
    .A1(\immu_1.page_table[1][9] ),
    .S(_1493_),
    .X(_1825_));
 sky130_fd_sc_hd__or2_1 _4321_ (.A(_1581_),
    .B(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__a31o_1 _4322_ (.A1(_1530_),
    .A2(_1824_),
    .A3(_1826_),
    .B1(_1553_),
    .X(_1827_));
 sky130_fd_sc_hd__o32a_1 _4323_ (.A1(_1457_),
    .A2(_1814_),
    .A3(_1818_),
    .B1(_1822_),
    .B2(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__a221oi_1 _4324_ (.A1(net107),
    .A2(_1810_),
    .B1(_1828_),
    .B2(_1441_),
    .C1(_0813_),
    .Y(_1829_));
 sky130_fd_sc_hd__nor2_2 _4325_ (.A(_1363_),
    .B(_1829_),
    .Y(_1830_));
 sky130_fd_sc_hd__a22o_4 _4326_ (.A1(_1569_),
    .A2(net244),
    .B1(_1805_),
    .B2(_1830_),
    .X(net678));
 sky130_fd_sc_hd__nand2_1 _4327_ (.A(net11),
    .B(\immu_0.high_addr_off[6] ),
    .Y(_1831_));
 sky130_fd_sc_hd__or2_1 _4328_ (.A(net11),
    .B(\immu_0.high_addr_off[6] ),
    .X(_1832_));
 sky130_fd_sc_hd__a21o_1 _4329_ (.A1(_1783_),
    .A2(_1785_),
    .B1(_1782_),
    .X(_1833_));
 sky130_fd_sc_hd__a21o_1 _4330_ (.A1(_1831_),
    .A2(_1832_),
    .B1(_1833_),
    .X(_1834_));
 sky130_fd_sc_hd__nand3_1 _4331_ (.A(_1831_),
    .B(_1832_),
    .C(_1833_),
    .Y(_1835_));
 sky130_fd_sc_hd__mux2_1 _4332_ (.A0(\immu_0.page_table[14][10] ),
    .A1(\immu_0.page_table[15][10] ),
    .S(_1480_),
    .X(_1836_));
 sky130_fd_sc_hd__nor2_1 _4333_ (.A(_1478_),
    .B(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hd__mux2_1 _4334_ (.A0(\immu_0.page_table[12][10] ),
    .A1(\immu_0.page_table[13][10] ),
    .S(_1408_),
    .X(_1838_));
 sky130_fd_sc_hd__o21ai_1 _4335_ (.A1(_1420_),
    .A2(_1838_),
    .B1(_1432_),
    .Y(_1839_));
 sky130_fd_sc_hd__mux2_1 _4336_ (.A0(\immu_0.page_table[8][10] ),
    .A1(\immu_0.page_table[9][10] ),
    .S(_1480_),
    .X(_1840_));
 sky130_fd_sc_hd__nor2_1 _4337_ (.A(_1570_),
    .B(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__mux2_1 _4338_ (.A0(\immu_0.page_table[10][10] ),
    .A1(\immu_0.page_table[11][10] ),
    .S(_1480_),
    .X(_1842_));
 sky130_fd_sc_hd__o21ai_1 _4339_ (.A1(_1478_),
    .A2(_1842_),
    .B1(_1535_),
    .Y(_1843_));
 sky130_fd_sc_hd__o221a_1 _4340_ (.A1(_1837_),
    .A2(_1839_),
    .B1(_1841_),
    .B2(_1843_),
    .C1(_1413_),
    .X(_1844_));
 sky130_fd_sc_hd__mux2_1 _4341_ (.A0(\immu_0.page_table[6][10] ),
    .A1(\immu_0.page_table[7][10] ),
    .S(_1425_),
    .X(_1845_));
 sky130_fd_sc_hd__or2_1 _4342_ (.A(_1424_),
    .B(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__mux2_1 _4343_ (.A0(\immu_0.page_table[4][10] ),
    .A1(\immu_0.page_table[5][10] ),
    .S(_1472_),
    .X(_1847_));
 sky130_fd_sc_hd__or2_1 _4344_ (.A(_1430_),
    .B(_1847_),
    .X(_1848_));
 sky130_fd_sc_hd__mux2_1 _4345_ (.A0(\immu_0.page_table[0][10] ),
    .A1(\immu_0.page_table[1][10] ),
    .S(_1425_),
    .X(_1849_));
 sky130_fd_sc_hd__mux2_1 _4346_ (.A0(\immu_0.page_table[2][10] ),
    .A1(\immu_0.page_table[3][10] ),
    .S(_1407_),
    .X(_1850_));
 sky130_fd_sc_hd__or2_1 _4347_ (.A(_1423_),
    .B(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__o211a_1 _4348_ (.A1(_1430_),
    .A2(_1849_),
    .B1(_1851_),
    .C1(_1416_),
    .X(_1852_));
 sky130_fd_sc_hd__a311o_1 _4349_ (.A1(_1432_),
    .A2(_1846_),
    .A3(_1848_),
    .B1(_1413_),
    .C1(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__and3b_1 _4350_ (.A_N(_1844_),
    .B(_1853_),
    .C(_1411_),
    .X(_1854_));
 sky130_fd_sc_hd__a311o_1 _4351_ (.A1(net2),
    .A2(_1834_),
    .A3(_1835_),
    .B1(_1854_),
    .C1(_1579_),
    .X(_1855_));
 sky130_fd_sc_hd__mux2_1 _4352_ (.A0(\immu_1.page_table[14][10] ),
    .A1(\immu_1.page_table[15][10] ),
    .S(_1524_),
    .X(_1856_));
 sky130_fd_sc_hd__or2_1 _4353_ (.A(_1523_),
    .B(_1856_),
    .X(_1857_));
 sky130_fd_sc_hd__mux2_1 _4354_ (.A0(\immu_1.page_table[12][10] ),
    .A1(\immu_1.page_table[13][10] ),
    .S(_1439_),
    .X(_1858_));
 sky130_fd_sc_hd__o21a_1 _4355_ (.A1(_1496_),
    .A2(_1858_),
    .B1(_1516_),
    .X(_1859_));
 sky130_fd_sc_hd__mux2_1 _4356_ (.A0(\immu_1.page_table[8][10] ),
    .A1(\immu_1.page_table[9][10] ),
    .S(_1439_),
    .X(_1860_));
 sky130_fd_sc_hd__or2_1 _4357_ (.A(_1496_),
    .B(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__mux2_1 _4358_ (.A0(\immu_1.page_table[10][10] ),
    .A1(\immu_1.page_table[11][10] ),
    .S(_1439_),
    .X(_1862_));
 sky130_fd_sc_hd__o21a_1 _4359_ (.A1(_1523_),
    .A2(_1862_),
    .B1(_1530_),
    .X(_1863_));
 sky130_fd_sc_hd__a221o_2 _4360_ (.A1(_1857_),
    .A2(_1859_),
    .B1(_1861_),
    .B2(_1863_),
    .C1(_1457_),
    .X(_1864_));
 sky130_fd_sc_hd__mux2_1 _4361_ (.A0(\immu_1.page_table[6][10] ),
    .A1(\immu_1.page_table[7][10] ),
    .S(_1524_),
    .X(_1865_));
 sky130_fd_sc_hd__or2_1 _4362_ (.A(_1523_),
    .B(_1865_),
    .X(_1866_));
 sky130_fd_sc_hd__mux2_1 _4363_ (.A0(\immu_1.page_table[4][10] ),
    .A1(\immu_1.page_table[5][10] ),
    .S(_1524_),
    .X(_1867_));
 sky130_fd_sc_hd__or2_1 _4364_ (.A(_1496_),
    .B(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__mux2_1 _4365_ (.A0(\immu_1.page_table[0][10] ),
    .A1(\immu_1.page_table[1][10] ),
    .S(_1439_),
    .X(_1869_));
 sky130_fd_sc_hd__mux2_1 _4366_ (.A0(\immu_1.page_table[2][10] ),
    .A1(\immu_1.page_table[3][10] ),
    .S(_1438_),
    .X(_1870_));
 sky130_fd_sc_hd__or2_1 _4367_ (.A(_1584_),
    .B(_1870_),
    .X(_1871_));
 sky130_fd_sc_hd__o211a_1 _4368_ (.A1(_1496_),
    .A2(_1869_),
    .B1(_1871_),
    .C1(_1530_),
    .X(_1872_));
 sky130_fd_sc_hd__a311o_1 _4369_ (.A1(_1516_),
    .A2(_1866_),
    .A3(_1868_),
    .B1(_1553_),
    .C1(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__nand2_1 _4370_ (.A(net116),
    .B(\immu_1.high_addr_off[6] ),
    .Y(_1874_));
 sky130_fd_sc_hd__or2_1 _4371_ (.A(net116),
    .B(\immu_1.high_addr_off[6] ),
    .X(_1875_));
 sky130_fd_sc_hd__and2_1 _4372_ (.A(_1807_),
    .B(_1809_),
    .X(_1876_));
 sky130_fd_sc_hd__a211o_1 _4373_ (.A1(_1874_),
    .A2(_1875_),
    .B1(_1876_),
    .C1(_1806_),
    .X(_1877_));
 sky130_fd_sc_hd__o211ai_1 _4374_ (.A1(_1806_),
    .A2(_1876_),
    .B1(_1875_),
    .C1(_1874_),
    .Y(_1878_));
 sky130_fd_sc_hd__and3_1 _4375_ (.A(net107),
    .B(_1877_),
    .C(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__a311o_2 _4376_ (.A1(_1441_),
    .A2(_1864_),
    .A3(_1873_),
    .B1(_1879_),
    .C1(_0813_),
    .X(_1880_));
 sky130_fd_sc_hd__and2_1 _4377_ (.A(\inner_wb_arbiter.o_sel_sig ),
    .B(net245),
    .X(_1881_));
 sky130_fd_sc_hd__a31o_4 _4378_ (.A1(net664),
    .A2(_1855_),
    .A3(_1880_),
    .B1(_1881_),
    .X(net679));
 sky130_fd_sc_hd__xor2_1 _4379_ (.A(net117),
    .B(\immu_1.high_addr_off[7] ),
    .X(_1882_));
 sky130_fd_sc_hd__a21oi_1 _4380_ (.A1(_1874_),
    .A2(_1878_),
    .B1(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__a31o_1 _4381_ (.A1(_1874_),
    .A2(_1878_),
    .A3(_1882_),
    .B1(_1440_),
    .X(_1884_));
 sky130_fd_sc_hd__nor3_4 _4382_ (.A(_0813_),
    .B(_1883_),
    .C(_1884_),
    .Y(_1885_));
 sky130_fd_sc_hd__xor2_1 _4383_ (.A(net12),
    .B(\immu_0.high_addr_off[7] ),
    .X(_1886_));
 sky130_fd_sc_hd__a21o_1 _4384_ (.A1(_1831_),
    .A2(_1835_),
    .B1(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__a31oi_1 _4385_ (.A1(_1831_),
    .A2(_1835_),
    .A3(_1886_),
    .B1(_1360_),
    .Y(_1888_));
 sky130_fd_sc_hd__a31o_1 _4386_ (.A1(net2),
    .A2(_1887_),
    .A3(_1888_),
    .B1(\inner_wb_arbiter.o_sel_sig ),
    .X(_1889_));
 sky130_fd_sc_hd__a2bb2o_4 _4387_ (.A1_N(_1885_),
    .A2_N(_1889_),
    .B1(_1569_),
    .B2(net246),
    .X(net680));
 sky130_fd_sc_hd__mux2_2 _4388_ (.A0(net329),
    .A1(net383),
    .S(_1390_),
    .X(_1890_));
 sky130_fd_sc_hd__mux2_4 _4389_ (.A0(net275),
    .A1(_1890_),
    .S(_0811_),
    .X(_1891_));
 sky130_fd_sc_hd__clkbuf_1 _4390_ (.A(_1891_),
    .X(net709));
 sky130_fd_sc_hd__mux2_2 _4391_ (.A0(net326),
    .A1(net380),
    .S(_0812_),
    .X(_1892_));
 sky130_fd_sc_hd__mux2_4 _4392_ (.A0(net272),
    .A1(_1892_),
    .S(_0811_),
    .X(_1893_));
 sky130_fd_sc_hd__clkbuf_1 _4393_ (.A(_1893_),
    .X(net706));
 sky130_fd_sc_hd__mux2_2 _4394_ (.A0(net327),
    .A1(net381),
    .S(_0812_),
    .X(_1894_));
 sky130_fd_sc_hd__mux2_4 _4395_ (.A0(net273),
    .A1(_1894_),
    .S(_0811_),
    .X(_1895_));
 sky130_fd_sc_hd__clkbuf_1 _4396_ (.A(_1895_),
    .X(net707));
 sky130_fd_sc_hd__inv_2 _4397_ (.A(net710),
    .Y(_1896_));
 sky130_fd_sc_hd__buf_6 _4398_ (.A(_1896_),
    .X(_1897_));
 sky130_fd_sc_hd__buf_6 _4399_ (.A(_1897_),
    .X(_1898_));
 sky130_fd_sc_hd__mux2_1 _4400_ (.A0(net325),
    .A1(net379),
    .S(\icache_arbiter.o_sel_sig ),
    .X(_1899_));
 sky130_fd_sc_hd__mux2_4 _4401_ (.A0(net255),
    .A1(_1899_),
    .S(_0811_),
    .X(_1900_));
 sky130_fd_sc_hd__and2_1 _4402_ (.A(_1898_),
    .B(_1900_),
    .X(_1901_));
 sky130_fd_sc_hd__clkbuf_1 _4403_ (.A(_1901_),
    .X(net689));
 sky130_fd_sc_hd__or2_1 _4404_ (.A(\icore_sregs.c1_disable ),
    .B(net384),
    .X(_1902_));
 sky130_fd_sc_hd__clkbuf_1 _4405_ (.A(_1902_),
    .X(net464));
 sky130_fd_sc_hd__and3_1 _4406_ (.A(net664),
    .B(_1579_),
    .C(net387),
    .X(_1903_));
 sky130_fd_sc_hd__clkbuf_1 _4407_ (.A(_1903_),
    .X(net645));
 sky130_fd_sc_hd__and3_1 _4408_ (.A(net664),
    .B(_1579_),
    .C(net388),
    .X(_1904_));
 sky130_fd_sc_hd__clkbuf_1 _4409_ (.A(_1904_),
    .X(net646));
 sky130_fd_sc_hd__and2_1 _4410_ (.A(net212),
    .B(_0835_),
    .X(_1905_));
 sky130_fd_sc_hd__clkbuf_2 _4411_ (.A(_1905_),
    .X(net468));
 sky130_fd_sc_hd__and2_1 _4412_ (.A(net213),
    .B(_0835_),
    .X(_1906_));
 sky130_fd_sc_hd__clkbuf_2 _4413_ (.A(_1906_),
    .X(net485));
 sky130_fd_sc_hd__and2_1 _4414_ (.A(_1373_),
    .B(net387),
    .X(_1907_));
 sky130_fd_sc_hd__clkbuf_1 _4415_ (.A(_1907_),
    .X(net567));
 sky130_fd_sc_hd__and2_1 _4416_ (.A(_1373_),
    .B(net388),
    .X(_1908_));
 sky130_fd_sc_hd__clkbuf_1 _4417_ (.A(_1908_),
    .X(net568));
 sky130_fd_sc_hd__and2_4 _4418_ (.A(_1373_),
    .B(net230),
    .X(_1909_));
 sky130_fd_sc_hd__clkbuf_1 _4419_ (.A(_1909_),
    .X(net663));
 sky130_fd_sc_hd__buf_4 _4420_ (.A(_1897_),
    .X(_1910_));
 sky130_fd_sc_hd__buf_8 _4421_ (.A(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__nand2_1 _4422_ (.A(net83),
    .B(net76),
    .Y(_1912_));
 sky130_fd_sc_hd__or2b_1 _4423_ (.A(net84),
    .B_N(net85),
    .X(_1913_));
 sky130_fd_sc_hd__or2_4 _4424_ (.A(_1912_),
    .B(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__or4_1 _4425_ (.A(net82),
    .B(net81),
    .C(net80),
    .D(net79),
    .X(_1915_));
 sky130_fd_sc_hd__or4b_1 _4426_ (.A(net78),
    .B(net77),
    .C(net91),
    .D_N(net90),
    .X(_1916_));
 sky130_fd_sc_hd__or2_1 _4427_ (.A(_1915_),
    .B(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__or4b_1 _4428_ (.A(net89),
    .B(net88),
    .C(net87),
    .D_N(net105),
    .X(_1918_));
 sky130_fd_sc_hd__or2_1 _4429_ (.A(net86),
    .B(_1918_),
    .X(_1919_));
 sky130_fd_sc_hd__or2_1 _4430_ (.A(net710),
    .B(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__or2_2 _4431_ (.A(_1917_),
    .B(_1920_),
    .X(_1921_));
 sky130_fd_sc_hd__buf_6 _4432_ (.A(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__or2_1 _4433_ (.A(_1914_),
    .B(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__buf_4 _4434_ (.A(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__inv_2 _4435_ (.A(net92),
    .Y(_1925_));
 sky130_fd_sc_hd__buf_4 _4436_ (.A(_1925_),
    .X(_1926_));
 sky130_fd_sc_hd__nor2_1 _4437_ (.A(_1926_),
    .B(_1923_),
    .Y(_1927_));
 sky130_fd_sc_hd__a31o_1 _4438_ (.A1(_1911_),
    .A2(\immu_0.page_table[11][0] ),
    .A3(_1924_),
    .B1(_1927_),
    .X(_0573_));
 sky130_fd_sc_hd__buf_6 _4439_ (.A(net96),
    .X(_1928_));
 sky130_fd_sc_hd__buf_4 _4440_ (.A(_1921_),
    .X(_1929_));
 sky130_fd_sc_hd__clkbuf_16 _4441_ (.A(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__nor2_4 _4442_ (.A(_1914_),
    .B(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__and2_1 _4443_ (.A(_1928_),
    .B(_1931_),
    .X(_1932_));
 sky130_fd_sc_hd__a31o_1 _4444_ (.A1(_1911_),
    .A2(\immu_0.page_table[11][1] ),
    .A3(_1924_),
    .B1(_1932_),
    .X(_0574_));
 sky130_fd_sc_hd__buf_6 _4445_ (.A(net97),
    .X(_1933_));
 sky130_fd_sc_hd__and2_1 _4446_ (.A(_1933_),
    .B(_1931_),
    .X(_1934_));
 sky130_fd_sc_hd__a31o_1 _4447_ (.A1(_1911_),
    .A2(\immu_0.page_table[11][2] ),
    .A3(_1924_),
    .B1(_1934_),
    .X(_0575_));
 sky130_fd_sc_hd__clkbuf_8 _4448_ (.A(net98),
    .X(_1935_));
 sky130_fd_sc_hd__and2_1 _4449_ (.A(_1935_),
    .B(_1931_),
    .X(_1936_));
 sky130_fd_sc_hd__a31o_1 _4450_ (.A1(_1911_),
    .A2(\immu_0.page_table[11][3] ),
    .A3(_1924_),
    .B1(_1936_),
    .X(_0576_));
 sky130_fd_sc_hd__buf_4 _4451_ (.A(net99),
    .X(_1937_));
 sky130_fd_sc_hd__and2_1 _4452_ (.A(_1937_),
    .B(_1931_),
    .X(_1938_));
 sky130_fd_sc_hd__a31o_1 _4453_ (.A1(_1911_),
    .A2(\immu_0.page_table[11][4] ),
    .A3(_1924_),
    .B1(_1938_),
    .X(_0577_));
 sky130_fd_sc_hd__buf_4 _4454_ (.A(_1898_),
    .X(_1939_));
 sky130_fd_sc_hd__buf_6 _4455_ (.A(net100),
    .X(_1940_));
 sky130_fd_sc_hd__and2_1 _4456_ (.A(_1940_),
    .B(_1931_),
    .X(_1941_));
 sky130_fd_sc_hd__a31o_1 _4457_ (.A1(_1939_),
    .A2(\immu_0.page_table[11][5] ),
    .A3(_1924_),
    .B1(_1941_),
    .X(_0578_));
 sky130_fd_sc_hd__buf_6 _4458_ (.A(net101),
    .X(_1942_));
 sky130_fd_sc_hd__and2_1 _4459_ (.A(_1942_),
    .B(_1931_),
    .X(_1943_));
 sky130_fd_sc_hd__a31o_1 _4460_ (.A1(_1939_),
    .A2(\immu_0.page_table[11][6] ),
    .A3(_1924_),
    .B1(_1943_),
    .X(_0579_));
 sky130_fd_sc_hd__buf_4 _4461_ (.A(net102),
    .X(_1944_));
 sky130_fd_sc_hd__and2_1 _4462_ (.A(_1944_),
    .B(_1931_),
    .X(_1945_));
 sky130_fd_sc_hd__a31o_1 _4463_ (.A1(_1939_),
    .A2(\immu_0.page_table[11][7] ),
    .A3(_1924_),
    .B1(_1945_),
    .X(_0580_));
 sky130_fd_sc_hd__buf_6 _4464_ (.A(net103),
    .X(_1946_));
 sky130_fd_sc_hd__and2_1 _4465_ (.A(_1946_),
    .B(_1931_),
    .X(_1947_));
 sky130_fd_sc_hd__a31o_1 _4466_ (.A1(_1939_),
    .A2(\immu_0.page_table[11][8] ),
    .A3(_1924_),
    .B1(_1947_),
    .X(_0581_));
 sky130_fd_sc_hd__buf_6 _4467_ (.A(net104),
    .X(_1948_));
 sky130_fd_sc_hd__and2_1 _4468_ (.A(_1948_),
    .B(_1931_),
    .X(_1949_));
 sky130_fd_sc_hd__a31o_1 _4469_ (.A1(_1939_),
    .A2(\immu_0.page_table[11][9] ),
    .A3(_1924_),
    .B1(_1949_),
    .X(_0582_));
 sky130_fd_sc_hd__buf_4 _4470_ (.A(net93),
    .X(_1950_));
 sky130_fd_sc_hd__and2_1 _4471_ (.A(_1950_),
    .B(_1931_),
    .X(_1951_));
 sky130_fd_sc_hd__a31o_1 _4472_ (.A1(_1939_),
    .A2(\immu_0.page_table[11][10] ),
    .A3(_1923_),
    .B1(_1951_),
    .X(_0583_));
 sky130_fd_sc_hd__or4_1 _4473_ (.A(net185),
    .B(net184),
    .C(net183),
    .D(net182),
    .X(_1952_));
 sky130_fd_sc_hd__or3_1 _4474_ (.A(net187),
    .B(net186),
    .C(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__or3b_4 _4475_ (.A(net195),
    .B(_1953_),
    .C_N(net196),
    .X(_1954_));
 sky130_fd_sc_hd__or4b_1 _4476_ (.A(net194),
    .B(net193),
    .C(net192),
    .D_N(net210),
    .X(_1955_));
 sky130_fd_sc_hd__or2_1 _4477_ (.A(net191),
    .B(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__or2_1 _4478_ (.A(net710),
    .B(_1956_),
    .X(_1957_));
 sky130_fd_sc_hd__or2_4 _4479_ (.A(_1954_),
    .B(_1957_),
    .X(_1958_));
 sky130_fd_sc_hd__or2b_1 _4480_ (.A(net181),
    .B_N(net188),
    .X(_1959_));
 sky130_fd_sc_hd__nand2_1 _4481_ (.A(net190),
    .B(net189),
    .Y(_1960_));
 sky130_fd_sc_hd__or2_2 _4482_ (.A(_1959_),
    .B(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__or2_1 _4483_ (.A(_1958_),
    .B(_1961_),
    .X(_1962_));
 sky130_fd_sc_hd__buf_2 _4484_ (.A(_1962_),
    .X(_1963_));
 sky130_fd_sc_hd__clkbuf_4 _4485_ (.A(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__inv_2 _4486_ (.A(net197),
    .Y(_1965_));
 sky130_fd_sc_hd__nor2_1 _4487_ (.A(_1965_),
    .B(_1963_),
    .Y(_1966_));
 sky130_fd_sc_hd__a31o_1 _4488_ (.A1(_1939_),
    .A2(\dmmu1.page_table[14][0] ),
    .A3(_1964_),
    .B1(_1966_),
    .X(_0584_));
 sky130_fd_sc_hd__buf_6 _4489_ (.A(net201),
    .X(_1967_));
 sky130_fd_sc_hd__clkbuf_4 _4490_ (.A(_1958_),
    .X(_1968_));
 sky130_fd_sc_hd__nor2_1 _4491_ (.A(_1968_),
    .B(_1961_),
    .Y(_1969_));
 sky130_fd_sc_hd__buf_2 _4492_ (.A(_1969_),
    .X(_1970_));
 sky130_fd_sc_hd__and2_1 _4493_ (.A(_1967_),
    .B(_1970_),
    .X(_1971_));
 sky130_fd_sc_hd__a31o_1 _4494_ (.A1(_1939_),
    .A2(\dmmu1.page_table[14][1] ),
    .A3(_1964_),
    .B1(_1971_),
    .X(_0585_));
 sky130_fd_sc_hd__buf_6 _4495_ (.A(net202),
    .X(_1972_));
 sky130_fd_sc_hd__and2_1 _4496_ (.A(_1972_),
    .B(_1970_),
    .X(_1973_));
 sky130_fd_sc_hd__a31o_1 _4497_ (.A1(_1939_),
    .A2(\dmmu1.page_table[14][2] ),
    .A3(_1964_),
    .B1(_1973_),
    .X(_0586_));
 sky130_fd_sc_hd__buf_6 _4498_ (.A(net203),
    .X(_1974_));
 sky130_fd_sc_hd__and2_1 _4499_ (.A(_1974_),
    .B(_1970_),
    .X(_1975_));
 sky130_fd_sc_hd__a31o_1 _4500_ (.A1(_1939_),
    .A2(\dmmu1.page_table[14][3] ),
    .A3(_1964_),
    .B1(_1975_),
    .X(_0587_));
 sky130_fd_sc_hd__buf_6 _4501_ (.A(_1898_),
    .X(_1976_));
 sky130_fd_sc_hd__buf_6 _4502_ (.A(net204),
    .X(_1977_));
 sky130_fd_sc_hd__and2_1 _4503_ (.A(_1977_),
    .B(_1970_),
    .X(_1978_));
 sky130_fd_sc_hd__a31o_1 _4504_ (.A1(_1976_),
    .A2(\dmmu1.page_table[14][4] ),
    .A3(_1964_),
    .B1(_1978_),
    .X(_0588_));
 sky130_fd_sc_hd__buf_6 _4505_ (.A(net205),
    .X(_1979_));
 sky130_fd_sc_hd__and2_1 _4506_ (.A(_1979_),
    .B(_1970_),
    .X(_1980_));
 sky130_fd_sc_hd__a31o_1 _4507_ (.A1(_1976_),
    .A2(\dmmu1.page_table[14][5] ),
    .A3(_1964_),
    .B1(_1980_),
    .X(_0589_));
 sky130_fd_sc_hd__buf_6 _4508_ (.A(net206),
    .X(_1981_));
 sky130_fd_sc_hd__and2_1 _4509_ (.A(_1981_),
    .B(_1970_),
    .X(_1982_));
 sky130_fd_sc_hd__a31o_1 _4510_ (.A1(_1976_),
    .A2(\dmmu1.page_table[14][6] ),
    .A3(_1964_),
    .B1(_1982_),
    .X(_0590_));
 sky130_fd_sc_hd__buf_6 _4511_ (.A(net207),
    .X(_1983_));
 sky130_fd_sc_hd__and2_1 _4512_ (.A(_1983_),
    .B(_1970_),
    .X(_1984_));
 sky130_fd_sc_hd__a31o_1 _4513_ (.A1(_1976_),
    .A2(\dmmu1.page_table[14][7] ),
    .A3(_1964_),
    .B1(_1984_),
    .X(_0591_));
 sky130_fd_sc_hd__buf_4 _4514_ (.A(net208),
    .X(_1985_));
 sky130_fd_sc_hd__and2_1 _4515_ (.A(_1985_),
    .B(_1970_),
    .X(_1986_));
 sky130_fd_sc_hd__a31o_1 _4516_ (.A1(_1976_),
    .A2(\dmmu1.page_table[14][8] ),
    .A3(_1964_),
    .B1(_1986_),
    .X(_0592_));
 sky130_fd_sc_hd__buf_4 _4517_ (.A(net209),
    .X(_1987_));
 sky130_fd_sc_hd__and2_1 _4518_ (.A(_1987_),
    .B(_1970_),
    .X(_1988_));
 sky130_fd_sc_hd__a31o_1 _4519_ (.A1(_1976_),
    .A2(\dmmu1.page_table[14][9] ),
    .A3(_1964_),
    .B1(_1988_),
    .X(_0593_));
 sky130_fd_sc_hd__buf_4 _4520_ (.A(net198),
    .X(_1989_));
 sky130_fd_sc_hd__and2_1 _4521_ (.A(_1989_),
    .B(_1970_),
    .X(_1990_));
 sky130_fd_sc_hd__a31o_1 _4522_ (.A1(_1976_),
    .A2(\dmmu1.page_table[14][10] ),
    .A3(_1963_),
    .B1(_1990_),
    .X(_0594_));
 sky130_fd_sc_hd__buf_2 _4523_ (.A(net199),
    .X(_1991_));
 sky130_fd_sc_hd__and2_1 _4524_ (.A(_1991_),
    .B(_1969_),
    .X(_1992_));
 sky130_fd_sc_hd__a31o_1 _4525_ (.A1(_1976_),
    .A2(\dmmu1.page_table[14][11] ),
    .A3(_1963_),
    .B1(_1992_),
    .X(_0595_));
 sky130_fd_sc_hd__buf_2 _4526_ (.A(net200),
    .X(_1993_));
 sky130_fd_sc_hd__and2_1 _4527_ (.A(_1993_),
    .B(_1969_),
    .X(_1994_));
 sky130_fd_sc_hd__a31o_1 _4528_ (.A1(_1976_),
    .A2(\dmmu1.page_table[14][12] ),
    .A3(_1963_),
    .B1(_1994_),
    .X(_0596_));
 sky130_fd_sc_hd__buf_6 _4529_ (.A(net197),
    .X(_1995_));
 sky130_fd_sc_hd__buf_6 _4530_ (.A(_1995_),
    .X(_1996_));
 sky130_fd_sc_hd__or3b_4 _4531_ (.A(_1953_),
    .B(net196),
    .C_N(net195),
    .X(_1997_));
 sky130_fd_sc_hd__or2_2 _4532_ (.A(_1957_),
    .B(_1997_),
    .X(_1998_));
 sky130_fd_sc_hd__clkbuf_4 _4533_ (.A(_1998_),
    .X(_1999_));
 sky130_fd_sc_hd__buf_4 _4534_ (.A(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__nor2_1 _4535_ (.A(_1961_),
    .B(_2000_),
    .Y(_2001_));
 sky130_fd_sc_hd__clkbuf_4 _4536_ (.A(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__or2_1 _4537_ (.A(_1961_),
    .B(_1998_),
    .X(_2003_));
 sky130_fd_sc_hd__clkbuf_4 _4538_ (.A(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__and3_1 _4539_ (.A(_1910_),
    .B(\immu_1.page_table[14][0] ),
    .C(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__a21o_1 _4540_ (.A1(_1996_),
    .A2(_2002_),
    .B1(_2005_),
    .X(_0597_));
 sky130_fd_sc_hd__buf_4 _4541_ (.A(_1967_),
    .X(_2006_));
 sky130_fd_sc_hd__and3_1 _4542_ (.A(_1910_),
    .B(\immu_1.page_table[14][1] ),
    .C(_2004_),
    .X(_2007_));
 sky130_fd_sc_hd__a21o_1 _4543_ (.A1(_2006_),
    .A2(_2002_),
    .B1(_2007_),
    .X(_0598_));
 sky130_fd_sc_hd__buf_6 _4544_ (.A(_1972_),
    .X(_2008_));
 sky130_fd_sc_hd__and3_1 _4545_ (.A(_1910_),
    .B(\immu_1.page_table[14][2] ),
    .C(_2004_),
    .X(_2009_));
 sky130_fd_sc_hd__a21o_1 _4546_ (.A1(_2008_),
    .A2(_2002_),
    .B1(_2009_),
    .X(_0599_));
 sky130_fd_sc_hd__buf_6 _4547_ (.A(_1974_),
    .X(_2010_));
 sky130_fd_sc_hd__and3_1 _4548_ (.A(_1910_),
    .B(\immu_1.page_table[14][3] ),
    .C(_2004_),
    .X(_2011_));
 sky130_fd_sc_hd__a21o_1 _4549_ (.A1(_2010_),
    .A2(_2002_),
    .B1(_2011_),
    .X(_0600_));
 sky130_fd_sc_hd__buf_6 _4550_ (.A(_1977_),
    .X(_2012_));
 sky130_fd_sc_hd__and3_1 _4551_ (.A(_1910_),
    .B(\immu_1.page_table[14][4] ),
    .C(_2004_),
    .X(_2013_));
 sky130_fd_sc_hd__a21o_1 _4552_ (.A1(_2012_),
    .A2(_2002_),
    .B1(_2013_),
    .X(_0601_));
 sky130_fd_sc_hd__buf_6 _4553_ (.A(_1979_),
    .X(_2014_));
 sky130_fd_sc_hd__and3_1 _4554_ (.A(_1910_),
    .B(\immu_1.page_table[14][5] ),
    .C(_2004_),
    .X(_2015_));
 sky130_fd_sc_hd__a21o_1 _4555_ (.A1(_2014_),
    .A2(_2002_),
    .B1(_2015_),
    .X(_0602_));
 sky130_fd_sc_hd__buf_6 _4556_ (.A(_1981_),
    .X(_2016_));
 sky130_fd_sc_hd__clkbuf_4 _4557_ (.A(_1897_),
    .X(_2017_));
 sky130_fd_sc_hd__and3_1 _4558_ (.A(_2017_),
    .B(\immu_1.page_table[14][6] ),
    .C(_2004_),
    .X(_2018_));
 sky130_fd_sc_hd__a21o_1 _4559_ (.A1(_2016_),
    .A2(_2002_),
    .B1(_2018_),
    .X(_0603_));
 sky130_fd_sc_hd__clkbuf_8 _4560_ (.A(_1983_),
    .X(_2019_));
 sky130_fd_sc_hd__and3_1 _4561_ (.A(_2017_),
    .B(\immu_1.page_table[14][7] ),
    .C(_2004_),
    .X(_2020_));
 sky130_fd_sc_hd__a21o_1 _4562_ (.A1(_2019_),
    .A2(_2002_),
    .B1(_2020_),
    .X(_0604_));
 sky130_fd_sc_hd__buf_4 _4563_ (.A(_1985_),
    .X(_2021_));
 sky130_fd_sc_hd__and3_1 _4564_ (.A(_2017_),
    .B(\immu_1.page_table[14][8] ),
    .C(_2004_),
    .X(_2022_));
 sky130_fd_sc_hd__a21o_1 _4565_ (.A1(_2021_),
    .A2(_2002_),
    .B1(_2022_),
    .X(_0605_));
 sky130_fd_sc_hd__clkbuf_8 _4566_ (.A(_1987_),
    .X(_2023_));
 sky130_fd_sc_hd__and3_1 _4567_ (.A(_2017_),
    .B(\immu_1.page_table[14][9] ),
    .C(_2004_),
    .X(_2024_));
 sky130_fd_sc_hd__a21o_1 _4568_ (.A1(_2023_),
    .A2(_2002_),
    .B1(_2024_),
    .X(_0606_));
 sky130_fd_sc_hd__buf_4 _4569_ (.A(_1989_),
    .X(_2025_));
 sky130_fd_sc_hd__and3_1 _4570_ (.A(_2017_),
    .B(\immu_1.page_table[14][10] ),
    .C(_2003_),
    .X(_2026_));
 sky130_fd_sc_hd__a21o_1 _4571_ (.A1(_2025_),
    .A2(_2001_),
    .B1(_2026_),
    .X(_0607_));
 sky130_fd_sc_hd__or2b_1 _4572_ (.A(net188),
    .B_N(net181),
    .X(_2027_));
 sky130_fd_sc_hd__or2_2 _4573_ (.A(_1960_),
    .B(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__nor2_1 _4574_ (.A(_2000_),
    .B(_2028_),
    .Y(_2029_));
 sky130_fd_sc_hd__clkbuf_4 _4575_ (.A(_2029_),
    .X(_2030_));
 sky130_fd_sc_hd__or2_1 _4576_ (.A(_1999_),
    .B(_2028_),
    .X(_2031_));
 sky130_fd_sc_hd__buf_2 _4577_ (.A(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__and3_1 _4578_ (.A(_2017_),
    .B(\immu_1.page_table[13][0] ),
    .C(_2032_),
    .X(_2033_));
 sky130_fd_sc_hd__a21o_1 _4579_ (.A1(_1996_),
    .A2(_2030_),
    .B1(_2033_),
    .X(_0608_));
 sky130_fd_sc_hd__and3_1 _4580_ (.A(_2017_),
    .B(\immu_1.page_table[13][1] ),
    .C(_2032_),
    .X(_2034_));
 sky130_fd_sc_hd__a21o_1 _4581_ (.A1(_2006_),
    .A2(_2030_),
    .B1(_2034_),
    .X(_0609_));
 sky130_fd_sc_hd__and3_1 _4582_ (.A(_2017_),
    .B(\immu_1.page_table[13][2] ),
    .C(_2032_),
    .X(_2035_));
 sky130_fd_sc_hd__a21o_1 _4583_ (.A1(_2008_),
    .A2(_2030_),
    .B1(_2035_),
    .X(_0610_));
 sky130_fd_sc_hd__and3_1 _4584_ (.A(_2017_),
    .B(\immu_1.page_table[13][3] ),
    .C(_2032_),
    .X(_2036_));
 sky130_fd_sc_hd__a21o_1 _4585_ (.A1(_2010_),
    .A2(_2030_),
    .B1(_2036_),
    .X(_0611_));
 sky130_fd_sc_hd__and3_1 _4586_ (.A(_2017_),
    .B(\immu_1.page_table[13][4] ),
    .C(_2032_),
    .X(_2037_));
 sky130_fd_sc_hd__a21o_1 _4587_ (.A1(_2012_),
    .A2(_2030_),
    .B1(_2037_),
    .X(_0612_));
 sky130_fd_sc_hd__buf_2 _4588_ (.A(_1897_),
    .X(_2038_));
 sky130_fd_sc_hd__and3_1 _4589_ (.A(_2038_),
    .B(\immu_1.page_table[13][5] ),
    .C(_2032_),
    .X(_2039_));
 sky130_fd_sc_hd__a21o_1 _4590_ (.A1(_2014_),
    .A2(_2030_),
    .B1(_2039_),
    .X(_0613_));
 sky130_fd_sc_hd__and3_1 _4591_ (.A(_2038_),
    .B(\immu_1.page_table[13][6] ),
    .C(_2032_),
    .X(_2040_));
 sky130_fd_sc_hd__a21o_1 _4592_ (.A1(_2016_),
    .A2(_2030_),
    .B1(_2040_),
    .X(_0614_));
 sky130_fd_sc_hd__and3_1 _4593_ (.A(_2038_),
    .B(\immu_1.page_table[13][7] ),
    .C(_2032_),
    .X(_2041_));
 sky130_fd_sc_hd__a21o_1 _4594_ (.A1(_2019_),
    .A2(_2030_),
    .B1(_2041_),
    .X(_0615_));
 sky130_fd_sc_hd__and3_1 _4595_ (.A(_2038_),
    .B(\immu_1.page_table[13][8] ),
    .C(_2032_),
    .X(_2042_));
 sky130_fd_sc_hd__a21o_1 _4596_ (.A1(_2021_),
    .A2(_2030_),
    .B1(_2042_),
    .X(_0616_));
 sky130_fd_sc_hd__and3_1 _4597_ (.A(_2038_),
    .B(\immu_1.page_table[13][9] ),
    .C(_2032_),
    .X(_2043_));
 sky130_fd_sc_hd__a21o_1 _4598_ (.A1(_2023_),
    .A2(_2030_),
    .B1(_2043_),
    .X(_0617_));
 sky130_fd_sc_hd__and3_1 _4599_ (.A(_2038_),
    .B(\immu_1.page_table[13][10] ),
    .C(_2031_),
    .X(_2044_));
 sky130_fd_sc_hd__a21o_1 _4600_ (.A1(_2025_),
    .A2(_2029_),
    .B1(_2044_),
    .X(_0618_));
 sky130_fd_sc_hd__or3_2 _4601_ (.A(net188),
    .B(net181),
    .C(_1960_),
    .X(_2045_));
 sky130_fd_sc_hd__nor2_1 _4602_ (.A(_2000_),
    .B(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__clkbuf_4 _4603_ (.A(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__or2_1 _4604_ (.A(_1999_),
    .B(_2045_),
    .X(_2048_));
 sky130_fd_sc_hd__buf_2 _4605_ (.A(_2048_),
    .X(_2049_));
 sky130_fd_sc_hd__and3_1 _4606_ (.A(_2038_),
    .B(\immu_1.page_table[12][0] ),
    .C(_2049_),
    .X(_2050_));
 sky130_fd_sc_hd__a21o_1 _4607_ (.A1(_1996_),
    .A2(_2047_),
    .B1(_2050_),
    .X(_0619_));
 sky130_fd_sc_hd__and3_1 _4608_ (.A(_2038_),
    .B(\immu_1.page_table[12][1] ),
    .C(_2049_),
    .X(_2051_));
 sky130_fd_sc_hd__a21o_1 _4609_ (.A1(_2006_),
    .A2(_2047_),
    .B1(_2051_),
    .X(_0620_));
 sky130_fd_sc_hd__and3_1 _4610_ (.A(_2038_),
    .B(\immu_1.page_table[12][2] ),
    .C(_2049_),
    .X(_2052_));
 sky130_fd_sc_hd__a21o_1 _4611_ (.A1(_2008_),
    .A2(_2047_),
    .B1(_2052_),
    .X(_0621_));
 sky130_fd_sc_hd__and3_1 _4612_ (.A(_2038_),
    .B(\immu_1.page_table[12][3] ),
    .C(_2049_),
    .X(_2053_));
 sky130_fd_sc_hd__a21o_1 _4613_ (.A1(_2010_),
    .A2(_2047_),
    .B1(_2053_),
    .X(_0622_));
 sky130_fd_sc_hd__buf_2 _4614_ (.A(_1897_),
    .X(_2054_));
 sky130_fd_sc_hd__and3_1 _4615_ (.A(_2054_),
    .B(\immu_1.page_table[12][4] ),
    .C(_2049_),
    .X(_2055_));
 sky130_fd_sc_hd__a21o_1 _4616_ (.A1(_2012_),
    .A2(_2047_),
    .B1(_2055_),
    .X(_0623_));
 sky130_fd_sc_hd__and3_1 _4617_ (.A(_2054_),
    .B(\immu_1.page_table[12][5] ),
    .C(_2049_),
    .X(_2056_));
 sky130_fd_sc_hd__a21o_1 _4618_ (.A1(_2014_),
    .A2(_2047_),
    .B1(_2056_),
    .X(_0624_));
 sky130_fd_sc_hd__and3_1 _4619_ (.A(_2054_),
    .B(\immu_1.page_table[12][6] ),
    .C(_2049_),
    .X(_2057_));
 sky130_fd_sc_hd__a21o_1 _4620_ (.A1(_2016_),
    .A2(_2047_),
    .B1(_2057_),
    .X(_0625_));
 sky130_fd_sc_hd__and3_1 _4621_ (.A(_2054_),
    .B(\immu_1.page_table[12][7] ),
    .C(_2049_),
    .X(_2058_));
 sky130_fd_sc_hd__a21o_1 _4622_ (.A1(_2019_),
    .A2(_2047_),
    .B1(_2058_),
    .X(_0626_));
 sky130_fd_sc_hd__and3_1 _4623_ (.A(_2054_),
    .B(\immu_1.page_table[12][8] ),
    .C(_2049_),
    .X(_2059_));
 sky130_fd_sc_hd__a21o_1 _4624_ (.A1(_2021_),
    .A2(_2047_),
    .B1(_2059_),
    .X(_0627_));
 sky130_fd_sc_hd__and3_1 _4625_ (.A(_2054_),
    .B(\immu_1.page_table[12][9] ),
    .C(_2049_),
    .X(_2060_));
 sky130_fd_sc_hd__a21o_1 _4626_ (.A1(_2023_),
    .A2(_2047_),
    .B1(_2060_),
    .X(_0628_));
 sky130_fd_sc_hd__and3_1 _4627_ (.A(_2054_),
    .B(\immu_1.page_table[12][10] ),
    .C(_2048_),
    .X(_2061_));
 sky130_fd_sc_hd__a21o_1 _4628_ (.A1(_2025_),
    .A2(_2046_),
    .B1(_2061_),
    .X(_0629_));
 sky130_fd_sc_hd__or2b_1 _4629_ (.A(net189),
    .B_N(net190),
    .X(_2062_));
 sky130_fd_sc_hd__nand2_1 _4630_ (.A(net188),
    .B(net181),
    .Y(_2063_));
 sky130_fd_sc_hd__or2_2 _4631_ (.A(_2062_),
    .B(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__nor2_1 _4632_ (.A(_2000_),
    .B(_2064_),
    .Y(_2065_));
 sky130_fd_sc_hd__clkbuf_4 _4633_ (.A(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__or2_1 _4634_ (.A(_1999_),
    .B(_2064_),
    .X(_2067_));
 sky130_fd_sc_hd__buf_2 _4635_ (.A(_2067_),
    .X(_2068_));
 sky130_fd_sc_hd__and3_1 _4636_ (.A(_2054_),
    .B(\immu_1.page_table[11][0] ),
    .C(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__a21o_1 _4637_ (.A1(_1996_),
    .A2(_2066_),
    .B1(_2069_),
    .X(_0630_));
 sky130_fd_sc_hd__and3_1 _4638_ (.A(_2054_),
    .B(\immu_1.page_table[11][1] ),
    .C(_2068_),
    .X(_2070_));
 sky130_fd_sc_hd__a21o_1 _4639_ (.A1(_2006_),
    .A2(_2066_),
    .B1(_2070_),
    .X(_0631_));
 sky130_fd_sc_hd__and3_1 _4640_ (.A(_2054_),
    .B(\immu_1.page_table[11][2] ),
    .C(_2068_),
    .X(_2071_));
 sky130_fd_sc_hd__a21o_1 _4641_ (.A1(_2008_),
    .A2(_2066_),
    .B1(_2071_),
    .X(_0632_));
 sky130_fd_sc_hd__buf_2 _4642_ (.A(_1897_),
    .X(_2072_));
 sky130_fd_sc_hd__and3_1 _4643_ (.A(_2072_),
    .B(\immu_1.page_table[11][3] ),
    .C(_2068_),
    .X(_2073_));
 sky130_fd_sc_hd__a21o_1 _4644_ (.A1(_2010_),
    .A2(_2066_),
    .B1(_2073_),
    .X(_0633_));
 sky130_fd_sc_hd__and3_1 _4645_ (.A(_2072_),
    .B(\immu_1.page_table[11][4] ),
    .C(_2068_),
    .X(_2074_));
 sky130_fd_sc_hd__a21o_1 _4646_ (.A1(_2012_),
    .A2(_2066_),
    .B1(_2074_),
    .X(_0634_));
 sky130_fd_sc_hd__and3_1 _4647_ (.A(_2072_),
    .B(\immu_1.page_table[11][5] ),
    .C(_2068_),
    .X(_2075_));
 sky130_fd_sc_hd__a21o_1 _4648_ (.A1(_2014_),
    .A2(_2066_),
    .B1(_2075_),
    .X(_0635_));
 sky130_fd_sc_hd__and3_1 _4649_ (.A(_2072_),
    .B(\immu_1.page_table[11][6] ),
    .C(_2068_),
    .X(_2076_));
 sky130_fd_sc_hd__a21o_1 _4650_ (.A1(_2016_),
    .A2(_2066_),
    .B1(_2076_),
    .X(_0636_));
 sky130_fd_sc_hd__and3_1 _4651_ (.A(_2072_),
    .B(\immu_1.page_table[11][7] ),
    .C(_2068_),
    .X(_2077_));
 sky130_fd_sc_hd__a21o_1 _4652_ (.A1(_2019_),
    .A2(_2066_),
    .B1(_2077_),
    .X(_0637_));
 sky130_fd_sc_hd__and3_1 _4653_ (.A(_2072_),
    .B(\immu_1.page_table[11][8] ),
    .C(_2068_),
    .X(_2078_));
 sky130_fd_sc_hd__a21o_1 _4654_ (.A1(_2021_),
    .A2(_2066_),
    .B1(_2078_),
    .X(_0638_));
 sky130_fd_sc_hd__and3_1 _4655_ (.A(_2072_),
    .B(\immu_1.page_table[11][9] ),
    .C(_2068_),
    .X(_2079_));
 sky130_fd_sc_hd__a21o_1 _4656_ (.A1(_2023_),
    .A2(_2066_),
    .B1(_2079_),
    .X(_0639_));
 sky130_fd_sc_hd__and3_1 _4657_ (.A(_2072_),
    .B(\immu_1.page_table[11][10] ),
    .C(_2067_),
    .X(_2080_));
 sky130_fd_sc_hd__a21o_1 _4658_ (.A1(_2025_),
    .A2(_2065_),
    .B1(_2080_),
    .X(_0640_));
 sky130_fd_sc_hd__or2_4 _4659_ (.A(_1959_),
    .B(_2062_),
    .X(_2081_));
 sky130_fd_sc_hd__nor2_1 _4660_ (.A(_2000_),
    .B(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__clkbuf_4 _4661_ (.A(_2082_),
    .X(_2083_));
 sky130_fd_sc_hd__clkbuf_4 _4662_ (.A(_1998_),
    .X(_2084_));
 sky130_fd_sc_hd__or2_1 _4663_ (.A(_2084_),
    .B(_2081_),
    .X(_2085_));
 sky130_fd_sc_hd__buf_2 _4664_ (.A(_2085_),
    .X(_2086_));
 sky130_fd_sc_hd__and3_1 _4665_ (.A(_2072_),
    .B(\immu_1.page_table[10][0] ),
    .C(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__a21o_1 _4666_ (.A1(_1996_),
    .A2(_2083_),
    .B1(_2087_),
    .X(_0641_));
 sky130_fd_sc_hd__and3_1 _4667_ (.A(_2072_),
    .B(\immu_1.page_table[10][1] ),
    .C(_2086_),
    .X(_2088_));
 sky130_fd_sc_hd__a21o_1 _4668_ (.A1(_2006_),
    .A2(_2083_),
    .B1(_2088_),
    .X(_0642_));
 sky130_fd_sc_hd__buf_2 _4669_ (.A(_1897_),
    .X(_2089_));
 sky130_fd_sc_hd__and3_1 _4670_ (.A(_2089_),
    .B(\immu_1.page_table[10][2] ),
    .C(_2086_),
    .X(_2090_));
 sky130_fd_sc_hd__a21o_1 _4671_ (.A1(_2008_),
    .A2(_2083_),
    .B1(_2090_),
    .X(_0643_));
 sky130_fd_sc_hd__and3_1 _4672_ (.A(_2089_),
    .B(\immu_1.page_table[10][3] ),
    .C(_2086_),
    .X(_2091_));
 sky130_fd_sc_hd__a21o_1 _4673_ (.A1(_2010_),
    .A2(_2083_),
    .B1(_2091_),
    .X(_0644_));
 sky130_fd_sc_hd__and3_1 _4674_ (.A(_2089_),
    .B(\immu_1.page_table[10][4] ),
    .C(_2086_),
    .X(_2092_));
 sky130_fd_sc_hd__a21o_1 _4675_ (.A1(_2012_),
    .A2(_2083_),
    .B1(_2092_),
    .X(_0645_));
 sky130_fd_sc_hd__and3_1 _4676_ (.A(_2089_),
    .B(\immu_1.page_table[10][5] ),
    .C(_2086_),
    .X(_2093_));
 sky130_fd_sc_hd__a21o_1 _4677_ (.A1(_2014_),
    .A2(_2083_),
    .B1(_2093_),
    .X(_0646_));
 sky130_fd_sc_hd__and3_1 _4678_ (.A(_2089_),
    .B(\immu_1.page_table[10][6] ),
    .C(_2086_),
    .X(_2094_));
 sky130_fd_sc_hd__a21o_1 _4679_ (.A1(_2016_),
    .A2(_2083_),
    .B1(_2094_),
    .X(_0647_));
 sky130_fd_sc_hd__and3_1 _4680_ (.A(_2089_),
    .B(\immu_1.page_table[10][7] ),
    .C(_2086_),
    .X(_2095_));
 sky130_fd_sc_hd__a21o_1 _4681_ (.A1(_2019_),
    .A2(_2083_),
    .B1(_2095_),
    .X(_0648_));
 sky130_fd_sc_hd__and3_1 _4682_ (.A(_2089_),
    .B(\immu_1.page_table[10][8] ),
    .C(_2086_),
    .X(_2096_));
 sky130_fd_sc_hd__a21o_1 _4683_ (.A1(_2021_),
    .A2(_2083_),
    .B1(_2096_),
    .X(_0649_));
 sky130_fd_sc_hd__and3_1 _4684_ (.A(_2089_),
    .B(\immu_1.page_table[10][9] ),
    .C(_2086_),
    .X(_2097_));
 sky130_fd_sc_hd__a21o_1 _4685_ (.A1(_2023_),
    .A2(_2083_),
    .B1(_2097_),
    .X(_0650_));
 sky130_fd_sc_hd__and3_1 _4686_ (.A(_2089_),
    .B(\immu_1.page_table[10][10] ),
    .C(_2085_),
    .X(_2098_));
 sky130_fd_sc_hd__a21o_1 _4687_ (.A1(_2025_),
    .A2(_2082_),
    .B1(_2098_),
    .X(_0651_));
 sky130_fd_sc_hd__or2_4 _4688_ (.A(_2027_),
    .B(_2062_),
    .X(_2099_));
 sky130_fd_sc_hd__nor2_1 _4689_ (.A(_2000_),
    .B(_2099_),
    .Y(_2100_));
 sky130_fd_sc_hd__clkbuf_4 _4690_ (.A(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__or2_1 _4691_ (.A(_2084_),
    .B(_2099_),
    .X(_2102_));
 sky130_fd_sc_hd__buf_2 _4692_ (.A(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__and3_1 _4693_ (.A(_2089_),
    .B(\immu_1.page_table[9][0] ),
    .C(_2103_),
    .X(_2104_));
 sky130_fd_sc_hd__a21o_1 _4694_ (.A1(_1996_),
    .A2(_2101_),
    .B1(_2104_),
    .X(_0652_));
 sky130_fd_sc_hd__buf_4 _4695_ (.A(_1896_),
    .X(_2105_));
 sky130_fd_sc_hd__buf_2 _4696_ (.A(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__and3_1 _4697_ (.A(_2106_),
    .B(\immu_1.page_table[9][1] ),
    .C(_2103_),
    .X(_2107_));
 sky130_fd_sc_hd__a21o_1 _4698_ (.A1(_2006_),
    .A2(_2101_),
    .B1(_2107_),
    .X(_0653_));
 sky130_fd_sc_hd__and3_1 _4699_ (.A(_2106_),
    .B(\immu_1.page_table[9][2] ),
    .C(_2103_),
    .X(_2108_));
 sky130_fd_sc_hd__a21o_1 _4700_ (.A1(_2008_),
    .A2(_2101_),
    .B1(_2108_),
    .X(_0654_));
 sky130_fd_sc_hd__and3_1 _4701_ (.A(_2106_),
    .B(\immu_1.page_table[9][3] ),
    .C(_2103_),
    .X(_2109_));
 sky130_fd_sc_hd__a21o_1 _4702_ (.A1(_2010_),
    .A2(_2101_),
    .B1(_2109_),
    .X(_0655_));
 sky130_fd_sc_hd__and3_1 _4703_ (.A(_2106_),
    .B(\immu_1.page_table[9][4] ),
    .C(_2103_),
    .X(_2110_));
 sky130_fd_sc_hd__a21o_1 _4704_ (.A1(_2012_),
    .A2(_2101_),
    .B1(_2110_),
    .X(_0656_));
 sky130_fd_sc_hd__and3_1 _4705_ (.A(_2106_),
    .B(\immu_1.page_table[9][5] ),
    .C(_2103_),
    .X(_2111_));
 sky130_fd_sc_hd__a21o_1 _4706_ (.A1(_2014_),
    .A2(_2101_),
    .B1(_2111_),
    .X(_0657_));
 sky130_fd_sc_hd__and3_1 _4707_ (.A(_2106_),
    .B(\immu_1.page_table[9][6] ),
    .C(_2103_),
    .X(_2112_));
 sky130_fd_sc_hd__a21o_1 _4708_ (.A1(_2016_),
    .A2(_2101_),
    .B1(_2112_),
    .X(_0658_));
 sky130_fd_sc_hd__and3_1 _4709_ (.A(_2106_),
    .B(\immu_1.page_table[9][7] ),
    .C(_2103_),
    .X(_2113_));
 sky130_fd_sc_hd__a21o_1 _4710_ (.A1(_2019_),
    .A2(_2101_),
    .B1(_2113_),
    .X(_0659_));
 sky130_fd_sc_hd__and3_1 _4711_ (.A(_2106_),
    .B(\immu_1.page_table[9][8] ),
    .C(_2103_),
    .X(_2114_));
 sky130_fd_sc_hd__a21o_1 _4712_ (.A1(_2021_),
    .A2(_2101_),
    .B1(_2114_),
    .X(_0660_));
 sky130_fd_sc_hd__and3_1 _4713_ (.A(_2106_),
    .B(\immu_1.page_table[9][9] ),
    .C(_2103_),
    .X(_2115_));
 sky130_fd_sc_hd__a21o_1 _4714_ (.A1(_2023_),
    .A2(_2101_),
    .B1(_2115_),
    .X(_0661_));
 sky130_fd_sc_hd__and3_1 _4715_ (.A(_2106_),
    .B(\immu_1.page_table[9][10] ),
    .C(_2102_),
    .X(_2116_));
 sky130_fd_sc_hd__a21o_1 _4716_ (.A1(_2025_),
    .A2(_2100_),
    .B1(_2116_),
    .X(_0662_));
 sky130_fd_sc_hd__or2b_1 _4717_ (.A(net190),
    .B_N(net189),
    .X(_2117_));
 sky130_fd_sc_hd__or2_4 _4718_ (.A(_1959_),
    .B(_2117_),
    .X(_2118_));
 sky130_fd_sc_hd__nor2_1 _4719_ (.A(_2000_),
    .B(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__clkbuf_4 _4720_ (.A(_2119_),
    .X(_2120_));
 sky130_fd_sc_hd__buf_2 _4721_ (.A(_2105_),
    .X(_2121_));
 sky130_fd_sc_hd__or2_1 _4722_ (.A(_2084_),
    .B(_2118_),
    .X(_2122_));
 sky130_fd_sc_hd__buf_2 _4723_ (.A(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__and3_1 _4724_ (.A(_2121_),
    .B(\immu_1.page_table[6][0] ),
    .C(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__a21o_1 _4725_ (.A1(_1996_),
    .A2(_2120_),
    .B1(_2124_),
    .X(_0663_));
 sky130_fd_sc_hd__and3_1 _4726_ (.A(_2121_),
    .B(\immu_1.page_table[6][1] ),
    .C(_2123_),
    .X(_2125_));
 sky130_fd_sc_hd__a21o_1 _4727_ (.A1(_2006_),
    .A2(_2120_),
    .B1(_2125_),
    .X(_0664_));
 sky130_fd_sc_hd__and3_1 _4728_ (.A(_2121_),
    .B(\immu_1.page_table[6][2] ),
    .C(_2123_),
    .X(_2126_));
 sky130_fd_sc_hd__a21o_1 _4729_ (.A1(_2008_),
    .A2(_2120_),
    .B1(_2126_),
    .X(_0665_));
 sky130_fd_sc_hd__and3_1 _4730_ (.A(_2121_),
    .B(\immu_1.page_table[6][3] ),
    .C(_2123_),
    .X(_2127_));
 sky130_fd_sc_hd__a21o_1 _4731_ (.A1(_2010_),
    .A2(_2120_),
    .B1(_2127_),
    .X(_0666_));
 sky130_fd_sc_hd__and3_1 _4732_ (.A(_2121_),
    .B(\immu_1.page_table[6][4] ),
    .C(_2123_),
    .X(_2128_));
 sky130_fd_sc_hd__a21o_1 _4733_ (.A1(_2012_),
    .A2(_2120_),
    .B1(_2128_),
    .X(_0667_));
 sky130_fd_sc_hd__and3_1 _4734_ (.A(_2121_),
    .B(\immu_1.page_table[6][5] ),
    .C(_2123_),
    .X(_2129_));
 sky130_fd_sc_hd__a21o_1 _4735_ (.A1(_2014_),
    .A2(_2120_),
    .B1(_2129_),
    .X(_0668_));
 sky130_fd_sc_hd__and3_1 _4736_ (.A(_2121_),
    .B(\immu_1.page_table[6][6] ),
    .C(_2123_),
    .X(_2130_));
 sky130_fd_sc_hd__a21o_1 _4737_ (.A1(_2016_),
    .A2(_2120_),
    .B1(_2130_),
    .X(_0669_));
 sky130_fd_sc_hd__and3_1 _4738_ (.A(_2121_),
    .B(\immu_1.page_table[6][7] ),
    .C(_2123_),
    .X(_2131_));
 sky130_fd_sc_hd__a21o_1 _4739_ (.A1(_2019_),
    .A2(_2120_),
    .B1(_2131_),
    .X(_0670_));
 sky130_fd_sc_hd__and3_1 _4740_ (.A(_2121_),
    .B(\immu_1.page_table[6][8] ),
    .C(_2123_),
    .X(_2132_));
 sky130_fd_sc_hd__a21o_1 _4741_ (.A1(_2021_),
    .A2(_2120_),
    .B1(_2132_),
    .X(_0671_));
 sky130_fd_sc_hd__and3_1 _4742_ (.A(_2121_),
    .B(\immu_1.page_table[6][9] ),
    .C(_2123_),
    .X(_2133_));
 sky130_fd_sc_hd__a21o_1 _4743_ (.A1(_2023_),
    .A2(_2120_),
    .B1(_2133_),
    .X(_0672_));
 sky130_fd_sc_hd__clkbuf_4 _4744_ (.A(_2105_),
    .X(_2134_));
 sky130_fd_sc_hd__and3_1 _4745_ (.A(_2134_),
    .B(\immu_1.page_table[6][10] ),
    .C(_2122_),
    .X(_2135_));
 sky130_fd_sc_hd__a21o_1 _4746_ (.A1(_2025_),
    .A2(_2119_),
    .B1(_2135_),
    .X(_0673_));
 sky130_fd_sc_hd__or2_4 _4747_ (.A(_2027_),
    .B(_2117_),
    .X(_2136_));
 sky130_fd_sc_hd__nor2_1 _4748_ (.A(_2000_),
    .B(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__clkbuf_4 _4749_ (.A(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__or2_1 _4750_ (.A(_2084_),
    .B(_2136_),
    .X(_2139_));
 sky130_fd_sc_hd__buf_2 _4751_ (.A(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__and3_1 _4752_ (.A(_2134_),
    .B(\immu_1.page_table[5][0] ),
    .C(_2140_),
    .X(_2141_));
 sky130_fd_sc_hd__a21o_1 _4753_ (.A1(_1996_),
    .A2(_2138_),
    .B1(_2141_),
    .X(_0674_));
 sky130_fd_sc_hd__and3_1 _4754_ (.A(_2134_),
    .B(\immu_1.page_table[5][1] ),
    .C(_2140_),
    .X(_2142_));
 sky130_fd_sc_hd__a21o_1 _4755_ (.A1(_2006_),
    .A2(_2138_),
    .B1(_2142_),
    .X(_0675_));
 sky130_fd_sc_hd__and3_1 _4756_ (.A(_2134_),
    .B(\immu_1.page_table[5][2] ),
    .C(_2140_),
    .X(_2143_));
 sky130_fd_sc_hd__a21o_1 _4757_ (.A1(_2008_),
    .A2(_2138_),
    .B1(_2143_),
    .X(_0676_));
 sky130_fd_sc_hd__and3_1 _4758_ (.A(_2134_),
    .B(\immu_1.page_table[5][3] ),
    .C(_2140_),
    .X(_2144_));
 sky130_fd_sc_hd__a21o_1 _4759_ (.A1(_2010_),
    .A2(_2138_),
    .B1(_2144_),
    .X(_0677_));
 sky130_fd_sc_hd__and3_1 _4760_ (.A(_2134_),
    .B(\immu_1.page_table[5][4] ),
    .C(_2140_),
    .X(_2145_));
 sky130_fd_sc_hd__a21o_1 _4761_ (.A1(_2012_),
    .A2(_2138_),
    .B1(_2145_),
    .X(_0678_));
 sky130_fd_sc_hd__and3_1 _4762_ (.A(_2134_),
    .B(\immu_1.page_table[5][5] ),
    .C(_2140_),
    .X(_2146_));
 sky130_fd_sc_hd__a21o_1 _4763_ (.A1(_2014_),
    .A2(_2138_),
    .B1(_2146_),
    .X(_0679_));
 sky130_fd_sc_hd__and3_1 _4764_ (.A(_2134_),
    .B(\immu_1.page_table[5][6] ),
    .C(_2140_),
    .X(_2147_));
 sky130_fd_sc_hd__a21o_1 _4765_ (.A1(_2016_),
    .A2(_2138_),
    .B1(_2147_),
    .X(_0680_));
 sky130_fd_sc_hd__and3_1 _4766_ (.A(_2134_),
    .B(\immu_1.page_table[5][7] ),
    .C(_2140_),
    .X(_2148_));
 sky130_fd_sc_hd__a21o_1 _4767_ (.A1(_2019_),
    .A2(_2138_),
    .B1(_2148_),
    .X(_0681_));
 sky130_fd_sc_hd__and3_1 _4768_ (.A(_2134_),
    .B(\immu_1.page_table[5][8] ),
    .C(_2140_),
    .X(_2149_));
 sky130_fd_sc_hd__a21o_1 _4769_ (.A1(_2021_),
    .A2(_2138_),
    .B1(_2149_),
    .X(_0682_));
 sky130_fd_sc_hd__buf_2 _4770_ (.A(_2105_),
    .X(_2150_));
 sky130_fd_sc_hd__and3_1 _4771_ (.A(_2150_),
    .B(\immu_1.page_table[5][9] ),
    .C(_2140_),
    .X(_2151_));
 sky130_fd_sc_hd__a21o_1 _4772_ (.A1(_2023_),
    .A2(_2138_),
    .B1(_2151_),
    .X(_0683_));
 sky130_fd_sc_hd__and3_1 _4773_ (.A(_2150_),
    .B(\immu_1.page_table[5][10] ),
    .C(_2139_),
    .X(_2152_));
 sky130_fd_sc_hd__a21o_1 _4774_ (.A1(_2025_),
    .A2(_2137_),
    .B1(_2152_),
    .X(_0684_));
 sky130_fd_sc_hd__or3_4 _4775_ (.A(net188),
    .B(net181),
    .C(_2117_),
    .X(_2153_));
 sky130_fd_sc_hd__nor2_1 _4776_ (.A(_2000_),
    .B(_2153_),
    .Y(_2154_));
 sky130_fd_sc_hd__clkbuf_4 _4777_ (.A(_2154_),
    .X(_2155_));
 sky130_fd_sc_hd__or2_1 _4778_ (.A(_2084_),
    .B(_2153_),
    .X(_2156_));
 sky130_fd_sc_hd__buf_2 _4779_ (.A(_2156_),
    .X(_2157_));
 sky130_fd_sc_hd__and3_1 _4780_ (.A(_2150_),
    .B(\immu_1.page_table[4][0] ),
    .C(_2157_),
    .X(_2158_));
 sky130_fd_sc_hd__a21o_1 _4781_ (.A1(_1996_),
    .A2(_2155_),
    .B1(_2158_),
    .X(_0685_));
 sky130_fd_sc_hd__and3_1 _4782_ (.A(_2150_),
    .B(\immu_1.page_table[4][1] ),
    .C(_2157_),
    .X(_2159_));
 sky130_fd_sc_hd__a21o_1 _4783_ (.A1(_2006_),
    .A2(_2155_),
    .B1(_2159_),
    .X(_0686_));
 sky130_fd_sc_hd__and3_1 _4784_ (.A(_2150_),
    .B(\immu_1.page_table[4][2] ),
    .C(_2157_),
    .X(_2160_));
 sky130_fd_sc_hd__a21o_1 _4785_ (.A1(_2008_),
    .A2(_2155_),
    .B1(_2160_),
    .X(_0687_));
 sky130_fd_sc_hd__and3_1 _4786_ (.A(_2150_),
    .B(\immu_1.page_table[4][3] ),
    .C(_2157_),
    .X(_2161_));
 sky130_fd_sc_hd__a21o_1 _4787_ (.A1(_2010_),
    .A2(_2155_),
    .B1(_2161_),
    .X(_0688_));
 sky130_fd_sc_hd__and3_1 _4788_ (.A(_2150_),
    .B(\immu_1.page_table[4][4] ),
    .C(_2157_),
    .X(_2162_));
 sky130_fd_sc_hd__a21o_1 _4789_ (.A1(_2012_),
    .A2(_2155_),
    .B1(_2162_),
    .X(_0689_));
 sky130_fd_sc_hd__and3_1 _4790_ (.A(_2150_),
    .B(\immu_1.page_table[4][5] ),
    .C(_2157_),
    .X(_2163_));
 sky130_fd_sc_hd__a21o_1 _4791_ (.A1(_2014_),
    .A2(_2155_),
    .B1(_2163_),
    .X(_0690_));
 sky130_fd_sc_hd__and3_1 _4792_ (.A(_2150_),
    .B(\immu_1.page_table[4][6] ),
    .C(_2157_),
    .X(_2164_));
 sky130_fd_sc_hd__a21o_1 _4793_ (.A1(_2016_),
    .A2(_2155_),
    .B1(_2164_),
    .X(_0691_));
 sky130_fd_sc_hd__and3_1 _4794_ (.A(_2150_),
    .B(\immu_1.page_table[4][7] ),
    .C(_2157_),
    .X(_2165_));
 sky130_fd_sc_hd__a21o_1 _4795_ (.A1(_2019_),
    .A2(_2155_),
    .B1(_2165_),
    .X(_0692_));
 sky130_fd_sc_hd__buf_2 _4796_ (.A(_2105_),
    .X(_2166_));
 sky130_fd_sc_hd__and3_1 _4797_ (.A(_2166_),
    .B(\immu_1.page_table[4][8] ),
    .C(_2157_),
    .X(_2167_));
 sky130_fd_sc_hd__a21o_1 _4798_ (.A1(_2021_),
    .A2(_2155_),
    .B1(_2167_),
    .X(_0693_));
 sky130_fd_sc_hd__and3_1 _4799_ (.A(_2166_),
    .B(\immu_1.page_table[4][9] ),
    .C(_2157_),
    .X(_2168_));
 sky130_fd_sc_hd__a21o_1 _4800_ (.A1(_2023_),
    .A2(_2155_),
    .B1(_2168_),
    .X(_0694_));
 sky130_fd_sc_hd__and3_1 _4801_ (.A(_2166_),
    .B(\immu_1.page_table[4][10] ),
    .C(_2156_),
    .X(_2169_));
 sky130_fd_sc_hd__a21o_1 _4802_ (.A1(_2025_),
    .A2(_2154_),
    .B1(_2169_),
    .X(_0695_));
 sky130_fd_sc_hd__or3_4 _4803_ (.A(net190),
    .B(net189),
    .C(_1959_),
    .X(_2170_));
 sky130_fd_sc_hd__nor2_1 _4804_ (.A(_2000_),
    .B(_2170_),
    .Y(_2171_));
 sky130_fd_sc_hd__clkbuf_4 _4805_ (.A(_2171_),
    .X(_2172_));
 sky130_fd_sc_hd__or2_1 _4806_ (.A(_2084_),
    .B(_2170_),
    .X(_2173_));
 sky130_fd_sc_hd__buf_2 _4807_ (.A(_2173_),
    .X(_2174_));
 sky130_fd_sc_hd__and3_1 _4808_ (.A(_2166_),
    .B(\immu_1.page_table[2][0] ),
    .C(_2174_),
    .X(_2175_));
 sky130_fd_sc_hd__a21o_1 _4809_ (.A1(_1996_),
    .A2(_2172_),
    .B1(_2175_),
    .X(_0696_));
 sky130_fd_sc_hd__and3_1 _4810_ (.A(_2166_),
    .B(\immu_1.page_table[2][1] ),
    .C(_2174_),
    .X(_2176_));
 sky130_fd_sc_hd__a21o_1 _4811_ (.A1(_2006_),
    .A2(_2172_),
    .B1(_2176_),
    .X(_0697_));
 sky130_fd_sc_hd__and3_1 _4812_ (.A(_2166_),
    .B(\immu_1.page_table[2][2] ),
    .C(_2174_),
    .X(_2177_));
 sky130_fd_sc_hd__a21o_1 _4813_ (.A1(_2008_),
    .A2(_2172_),
    .B1(_2177_),
    .X(_0698_));
 sky130_fd_sc_hd__and3_1 _4814_ (.A(_2166_),
    .B(\immu_1.page_table[2][3] ),
    .C(_2174_),
    .X(_2178_));
 sky130_fd_sc_hd__a21o_1 _4815_ (.A1(_2010_),
    .A2(_2172_),
    .B1(_2178_),
    .X(_0699_));
 sky130_fd_sc_hd__and3_1 _4816_ (.A(_2166_),
    .B(\immu_1.page_table[2][4] ),
    .C(_2174_),
    .X(_2179_));
 sky130_fd_sc_hd__a21o_1 _4817_ (.A1(_2012_),
    .A2(_2172_),
    .B1(_2179_),
    .X(_0700_));
 sky130_fd_sc_hd__and3_1 _4818_ (.A(_2166_),
    .B(\immu_1.page_table[2][5] ),
    .C(_2174_),
    .X(_2180_));
 sky130_fd_sc_hd__a21o_1 _4819_ (.A1(_2014_),
    .A2(_2172_),
    .B1(_2180_),
    .X(_0701_));
 sky130_fd_sc_hd__and3_1 _4820_ (.A(_2166_),
    .B(\immu_1.page_table[2][6] ),
    .C(_2174_),
    .X(_2181_));
 sky130_fd_sc_hd__a21o_1 _4821_ (.A1(_2016_),
    .A2(_2172_),
    .B1(_2181_),
    .X(_0702_));
 sky130_fd_sc_hd__buf_2 _4822_ (.A(_2105_),
    .X(_2182_));
 sky130_fd_sc_hd__and3_1 _4823_ (.A(_2182_),
    .B(\immu_1.page_table[2][7] ),
    .C(_2174_),
    .X(_2183_));
 sky130_fd_sc_hd__a21o_1 _4824_ (.A1(_2019_),
    .A2(_2172_),
    .B1(_2183_),
    .X(_0703_));
 sky130_fd_sc_hd__and3_1 _4825_ (.A(_2182_),
    .B(\immu_1.page_table[2][8] ),
    .C(_2174_),
    .X(_2184_));
 sky130_fd_sc_hd__a21o_1 _4826_ (.A1(_2021_),
    .A2(_2172_),
    .B1(_2184_),
    .X(_0704_));
 sky130_fd_sc_hd__and3_1 _4827_ (.A(_2182_),
    .B(\immu_1.page_table[2][9] ),
    .C(_2174_),
    .X(_2185_));
 sky130_fd_sc_hd__a21o_1 _4828_ (.A1(_2023_),
    .A2(_2172_),
    .B1(_2185_),
    .X(_0705_));
 sky130_fd_sc_hd__and3_1 _4829_ (.A(_2182_),
    .B(\immu_1.page_table[2][10] ),
    .C(_2173_),
    .X(_2186_));
 sky130_fd_sc_hd__a21o_1 _4830_ (.A1(_2025_),
    .A2(_2171_),
    .B1(_2186_),
    .X(_0706_));
 sky130_fd_sc_hd__or3_2 _4831_ (.A(net190),
    .B(net189),
    .C(_2027_),
    .X(_2187_));
 sky130_fd_sc_hd__or2_1 _4832_ (.A(_1999_),
    .B(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__buf_4 _4833_ (.A(_2188_),
    .X(_2189_));
 sky130_fd_sc_hd__buf_4 _4834_ (.A(_1896_),
    .X(_2190_));
 sky130_fd_sc_hd__nand2_1 _4835_ (.A(_2190_),
    .B(_2188_),
    .Y(_2191_));
 sky130_fd_sc_hd__clkbuf_4 _4836_ (.A(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__o22a_1 _4837_ (.A1(_1995_),
    .A2(_2189_),
    .B1(_2192_),
    .B2(\immu_1.page_table[1][0] ),
    .X(_0707_));
 sky130_fd_sc_hd__o22a_1 _4838_ (.A1(_1967_),
    .A2(_2189_),
    .B1(_2192_),
    .B2(\immu_1.page_table[1][1] ),
    .X(_0708_));
 sky130_fd_sc_hd__o22a_1 _4839_ (.A1(_1972_),
    .A2(_2189_),
    .B1(_2192_),
    .B2(\immu_1.page_table[1][2] ),
    .X(_0709_));
 sky130_fd_sc_hd__o22a_1 _4840_ (.A1(_1974_),
    .A2(_2189_),
    .B1(_2192_),
    .B2(\immu_1.page_table[1][3] ),
    .X(_0710_));
 sky130_fd_sc_hd__o22a_1 _4841_ (.A1(_1977_),
    .A2(_2189_),
    .B1(_2192_),
    .B2(\immu_1.page_table[1][4] ),
    .X(_0711_));
 sky130_fd_sc_hd__o22a_1 _4842_ (.A1(_1979_),
    .A2(_2189_),
    .B1(_2192_),
    .B2(\immu_1.page_table[1][5] ),
    .X(_0712_));
 sky130_fd_sc_hd__o22a_1 _4843_ (.A1(_1981_),
    .A2(_2189_),
    .B1(_2192_),
    .B2(\immu_1.page_table[1][6] ),
    .X(_0713_));
 sky130_fd_sc_hd__o22a_1 _4844_ (.A1(_1983_),
    .A2(_2189_),
    .B1(_2192_),
    .B2(\immu_1.page_table[1][7] ),
    .X(_0714_));
 sky130_fd_sc_hd__o22a_1 _4845_ (.A1(_1985_),
    .A2(_2189_),
    .B1(_2192_),
    .B2(\immu_1.page_table[1][8] ),
    .X(_0715_));
 sky130_fd_sc_hd__o22a_1 _4846_ (.A1(_1987_),
    .A2(_2189_),
    .B1(_2192_),
    .B2(\immu_1.page_table[1][9] ),
    .X(_0716_));
 sky130_fd_sc_hd__o22a_1 _4847_ (.A1(_1989_),
    .A2(_2188_),
    .B1(_2191_),
    .B2(\immu_1.page_table[1][10] ),
    .X(_0717_));
 sky130_fd_sc_hd__or3_4 _4848_ (.A(net190),
    .B(net189),
    .C(_2063_),
    .X(_2193_));
 sky130_fd_sc_hd__nor2_1 _4849_ (.A(_1999_),
    .B(_2193_),
    .Y(_2194_));
 sky130_fd_sc_hd__clkbuf_4 _4850_ (.A(_2194_),
    .X(_2195_));
 sky130_fd_sc_hd__or2_1 _4851_ (.A(_2084_),
    .B(_2193_),
    .X(_2196_));
 sky130_fd_sc_hd__buf_2 _4852_ (.A(_2196_),
    .X(_2197_));
 sky130_fd_sc_hd__and3_1 _4853_ (.A(_2182_),
    .B(\immu_1.page_table[3][0] ),
    .C(_2197_),
    .X(_2198_));
 sky130_fd_sc_hd__a21o_1 _4854_ (.A1(_1995_),
    .A2(_2195_),
    .B1(_2198_),
    .X(_0718_));
 sky130_fd_sc_hd__and3_1 _4855_ (.A(_2182_),
    .B(\immu_1.page_table[3][1] ),
    .C(_2197_),
    .X(_2199_));
 sky130_fd_sc_hd__a21o_1 _4856_ (.A1(_1967_),
    .A2(_2195_),
    .B1(_2199_),
    .X(_0719_));
 sky130_fd_sc_hd__and3_1 _4857_ (.A(_2182_),
    .B(\immu_1.page_table[3][2] ),
    .C(_2197_),
    .X(_2200_));
 sky130_fd_sc_hd__a21o_1 _4858_ (.A1(_1972_),
    .A2(_2195_),
    .B1(_2200_),
    .X(_0720_));
 sky130_fd_sc_hd__and3_1 _4859_ (.A(_2182_),
    .B(\immu_1.page_table[3][3] ),
    .C(_2197_),
    .X(_2201_));
 sky130_fd_sc_hd__a21o_1 _4860_ (.A1(_1974_),
    .A2(_2195_),
    .B1(_2201_),
    .X(_0721_));
 sky130_fd_sc_hd__and3_1 _4861_ (.A(_2182_),
    .B(\immu_1.page_table[3][4] ),
    .C(_2197_),
    .X(_2202_));
 sky130_fd_sc_hd__a21o_1 _4862_ (.A1(_1977_),
    .A2(_2195_),
    .B1(_2202_),
    .X(_0722_));
 sky130_fd_sc_hd__and3_1 _4863_ (.A(_2182_),
    .B(\immu_1.page_table[3][5] ),
    .C(_2197_),
    .X(_2203_));
 sky130_fd_sc_hd__a21o_1 _4864_ (.A1(_1979_),
    .A2(_2195_),
    .B1(_2203_),
    .X(_0723_));
 sky130_fd_sc_hd__buf_4 _4865_ (.A(_2105_),
    .X(_2204_));
 sky130_fd_sc_hd__and3_1 _4866_ (.A(_2204_),
    .B(\immu_1.page_table[3][6] ),
    .C(_2197_),
    .X(_2205_));
 sky130_fd_sc_hd__a21o_1 _4867_ (.A1(_1981_),
    .A2(_2195_),
    .B1(_2205_),
    .X(_0724_));
 sky130_fd_sc_hd__and3_1 _4868_ (.A(_2204_),
    .B(\immu_1.page_table[3][7] ),
    .C(_2197_),
    .X(_2206_));
 sky130_fd_sc_hd__a21o_1 _4869_ (.A1(_1983_),
    .A2(_2195_),
    .B1(_2206_),
    .X(_0725_));
 sky130_fd_sc_hd__and3_1 _4870_ (.A(_2204_),
    .B(\immu_1.page_table[3][8] ),
    .C(_2197_),
    .X(_2207_));
 sky130_fd_sc_hd__a21o_1 _4871_ (.A1(_1985_),
    .A2(_2195_),
    .B1(_2207_),
    .X(_0726_));
 sky130_fd_sc_hd__and3_1 _4872_ (.A(_2204_),
    .B(\immu_1.page_table[3][9] ),
    .C(_2197_),
    .X(_2208_));
 sky130_fd_sc_hd__a21o_1 _4873_ (.A1(_1987_),
    .A2(_2195_),
    .B1(_2208_),
    .X(_0727_));
 sky130_fd_sc_hd__and3_1 _4874_ (.A(_2204_),
    .B(\immu_1.page_table[3][10] ),
    .C(_2196_),
    .X(_2209_));
 sky130_fd_sc_hd__a21o_1 _4875_ (.A1(_1989_),
    .A2(_2194_),
    .B1(_2209_),
    .X(_0728_));
 sky130_fd_sc_hd__buf_6 _4876_ (.A(net92),
    .X(_2210_));
 sky130_fd_sc_hd__buf_4 _4877_ (.A(_2210_),
    .X(_2211_));
 sky130_fd_sc_hd__or4_4 _4878_ (.A(net83),
    .B(net76),
    .C(net85),
    .D(net84),
    .X(_2212_));
 sky130_fd_sc_hd__or2_1 _4879_ (.A(net90),
    .B(_1915_),
    .X(_2213_));
 sky130_fd_sc_hd__or4b_2 _4880_ (.A(net78),
    .B(_2213_),
    .C(net77),
    .D_N(net91),
    .X(_2214_));
 sky130_fd_sc_hd__or2_2 _4881_ (.A(_1920_),
    .B(_2214_),
    .X(_2215_));
 sky130_fd_sc_hd__buf_4 _4882_ (.A(_2215_),
    .X(_2216_));
 sky130_fd_sc_hd__buf_4 _4883_ (.A(_2216_),
    .X(_2217_));
 sky130_fd_sc_hd__nor2_1 _4884_ (.A(_2212_),
    .B(_2217_),
    .Y(_2218_));
 sky130_fd_sc_hd__buf_4 _4885_ (.A(_2218_),
    .X(_2219_));
 sky130_fd_sc_hd__or2_1 _4886_ (.A(_2212_),
    .B(_2215_),
    .X(_2220_));
 sky130_fd_sc_hd__clkbuf_4 _4887_ (.A(_2220_),
    .X(_2221_));
 sky130_fd_sc_hd__and3_1 _4888_ (.A(_2204_),
    .B(\dmmu0.page_table[0][0] ),
    .C(_2221_),
    .X(_2222_));
 sky130_fd_sc_hd__a21o_1 _4889_ (.A1(_2211_),
    .A2(_2219_),
    .B1(_2222_),
    .X(_0729_));
 sky130_fd_sc_hd__buf_8 _4890_ (.A(net96),
    .X(_2223_));
 sky130_fd_sc_hd__buf_4 _4891_ (.A(_2223_),
    .X(_2224_));
 sky130_fd_sc_hd__and3_1 _4892_ (.A(_2204_),
    .B(\dmmu0.page_table[0][1] ),
    .C(_2221_),
    .X(_2225_));
 sky130_fd_sc_hd__a21o_1 _4893_ (.A1(_2224_),
    .A2(_2219_),
    .B1(_2225_),
    .X(_0730_));
 sky130_fd_sc_hd__buf_4 _4894_ (.A(net97),
    .X(_2226_));
 sky130_fd_sc_hd__clkbuf_4 _4895_ (.A(_2226_),
    .X(_2227_));
 sky130_fd_sc_hd__and3_1 _4896_ (.A(_2204_),
    .B(\dmmu0.page_table[0][2] ),
    .C(_2221_),
    .X(_2228_));
 sky130_fd_sc_hd__a21o_1 _4897_ (.A1(_2227_),
    .A2(_2219_),
    .B1(_2228_),
    .X(_0731_));
 sky130_fd_sc_hd__buf_6 _4898_ (.A(net98),
    .X(_2229_));
 sky130_fd_sc_hd__buf_4 _4899_ (.A(_2229_),
    .X(_2230_));
 sky130_fd_sc_hd__and3_1 _4900_ (.A(_2204_),
    .B(\dmmu0.page_table[0][3] ),
    .C(_2221_),
    .X(_2231_));
 sky130_fd_sc_hd__a21o_1 _4901_ (.A1(_2230_),
    .A2(_2219_),
    .B1(_2231_),
    .X(_0732_));
 sky130_fd_sc_hd__buf_4 _4902_ (.A(net99),
    .X(_2232_));
 sky130_fd_sc_hd__buf_4 _4903_ (.A(_2232_),
    .X(_2233_));
 sky130_fd_sc_hd__and3_1 _4904_ (.A(_2204_),
    .B(\dmmu0.page_table[0][4] ),
    .C(_2221_),
    .X(_2234_));
 sky130_fd_sc_hd__a21o_1 _4905_ (.A1(_2233_),
    .A2(_2219_),
    .B1(_2234_),
    .X(_0733_));
 sky130_fd_sc_hd__buf_6 _4906_ (.A(net100),
    .X(_2235_));
 sky130_fd_sc_hd__buf_4 _4907_ (.A(_2235_),
    .X(_2236_));
 sky130_fd_sc_hd__clkbuf_4 _4908_ (.A(_2105_),
    .X(_2237_));
 sky130_fd_sc_hd__and3_1 _4909_ (.A(_2237_),
    .B(\dmmu0.page_table[0][5] ),
    .C(_2221_),
    .X(_2238_));
 sky130_fd_sc_hd__a21o_1 _4910_ (.A1(_2236_),
    .A2(_2219_),
    .B1(_2238_),
    .X(_0734_));
 sky130_fd_sc_hd__buf_6 _4911_ (.A(net101),
    .X(_2239_));
 sky130_fd_sc_hd__buf_4 _4912_ (.A(_2239_),
    .X(_2240_));
 sky130_fd_sc_hd__and3_1 _4913_ (.A(_2237_),
    .B(\dmmu0.page_table[0][6] ),
    .C(_2221_),
    .X(_2241_));
 sky130_fd_sc_hd__a21o_1 _4914_ (.A1(_2240_),
    .A2(_2219_),
    .B1(_2241_),
    .X(_0735_));
 sky130_fd_sc_hd__buf_6 _4915_ (.A(net102),
    .X(_2242_));
 sky130_fd_sc_hd__buf_4 _4916_ (.A(_2242_),
    .X(_2243_));
 sky130_fd_sc_hd__and3_1 _4917_ (.A(_2237_),
    .B(\dmmu0.page_table[0][7] ),
    .C(_2221_),
    .X(_2244_));
 sky130_fd_sc_hd__a21o_1 _4918_ (.A1(_2243_),
    .A2(_2219_),
    .B1(_2244_),
    .X(_0736_));
 sky130_fd_sc_hd__buf_6 _4919_ (.A(_1946_),
    .X(_2245_));
 sky130_fd_sc_hd__and3_1 _4920_ (.A(_2237_),
    .B(\dmmu0.page_table[0][8] ),
    .C(_2221_),
    .X(_2246_));
 sky130_fd_sc_hd__a21o_1 _4921_ (.A1(_2245_),
    .A2(_2219_),
    .B1(_2246_),
    .X(_0737_));
 sky130_fd_sc_hd__buf_4 _4922_ (.A(_1948_),
    .X(_2247_));
 sky130_fd_sc_hd__and3_1 _4923_ (.A(_2237_),
    .B(\dmmu0.page_table[0][9] ),
    .C(_2221_),
    .X(_2248_));
 sky130_fd_sc_hd__a21o_1 _4924_ (.A1(_2247_),
    .A2(_2219_),
    .B1(_2248_),
    .X(_0738_));
 sky130_fd_sc_hd__buf_4 _4925_ (.A(_1950_),
    .X(_2249_));
 sky130_fd_sc_hd__and3_1 _4926_ (.A(_2237_),
    .B(\dmmu0.page_table[0][10] ),
    .C(_2220_),
    .X(_2250_));
 sky130_fd_sc_hd__a21o_1 _4927_ (.A1(_2249_),
    .A2(_2218_),
    .B1(_2250_),
    .X(_0739_));
 sky130_fd_sc_hd__buf_4 _4928_ (.A(net94),
    .X(_2251_));
 sky130_fd_sc_hd__and3_1 _4929_ (.A(_2237_),
    .B(\dmmu0.page_table[0][11] ),
    .C(_2220_),
    .X(_2252_));
 sky130_fd_sc_hd__a21o_1 _4930_ (.A1(_2251_),
    .A2(_2218_),
    .B1(_2252_),
    .X(_0740_));
 sky130_fd_sc_hd__buf_4 _4931_ (.A(net95),
    .X(_2253_));
 sky130_fd_sc_hd__and3_1 _4932_ (.A(_2237_),
    .B(\dmmu0.page_table[0][12] ),
    .C(_2220_),
    .X(_2254_));
 sky130_fd_sc_hd__a21o_1 _4933_ (.A1(_2253_),
    .A2(_2218_),
    .B1(_2254_),
    .X(_0741_));
 sky130_fd_sc_hd__or2_2 _4934_ (.A(_2063_),
    .B(_2117_),
    .X(_2255_));
 sky130_fd_sc_hd__nor2_1 _4935_ (.A(_1999_),
    .B(_2255_),
    .Y(_2256_));
 sky130_fd_sc_hd__clkbuf_4 _4936_ (.A(_2256_),
    .X(_2257_));
 sky130_fd_sc_hd__or2_1 _4937_ (.A(_2084_),
    .B(_2255_),
    .X(_2258_));
 sky130_fd_sc_hd__buf_2 _4938_ (.A(_2258_),
    .X(_2259_));
 sky130_fd_sc_hd__and3_1 _4939_ (.A(_2237_),
    .B(\immu_1.page_table[7][0] ),
    .C(_2259_),
    .X(_2260_));
 sky130_fd_sc_hd__a21o_1 _4940_ (.A1(_1995_),
    .A2(_2257_),
    .B1(_2260_),
    .X(_0742_));
 sky130_fd_sc_hd__and3_1 _4941_ (.A(_2237_),
    .B(\immu_1.page_table[7][1] ),
    .C(_2259_),
    .X(_2261_));
 sky130_fd_sc_hd__a21o_1 _4942_ (.A1(_1967_),
    .A2(_2257_),
    .B1(_2261_),
    .X(_0743_));
 sky130_fd_sc_hd__clkbuf_4 _4943_ (.A(_2105_),
    .X(_2262_));
 sky130_fd_sc_hd__and3_1 _4944_ (.A(_2262_),
    .B(\immu_1.page_table[7][2] ),
    .C(_2259_),
    .X(_2263_));
 sky130_fd_sc_hd__a21o_1 _4945_ (.A1(_1972_),
    .A2(_2257_),
    .B1(_2263_),
    .X(_0744_));
 sky130_fd_sc_hd__and3_1 _4946_ (.A(_2262_),
    .B(\immu_1.page_table[7][3] ),
    .C(_2259_),
    .X(_2264_));
 sky130_fd_sc_hd__a21o_1 _4947_ (.A1(_1974_),
    .A2(_2257_),
    .B1(_2264_),
    .X(_0745_));
 sky130_fd_sc_hd__and3_1 _4948_ (.A(_2262_),
    .B(\immu_1.page_table[7][4] ),
    .C(_2259_),
    .X(_2265_));
 sky130_fd_sc_hd__a21o_1 _4949_ (.A1(_1977_),
    .A2(_2257_),
    .B1(_2265_),
    .X(_0746_));
 sky130_fd_sc_hd__and3_1 _4950_ (.A(_2262_),
    .B(\immu_1.page_table[7][5] ),
    .C(_2259_),
    .X(_2266_));
 sky130_fd_sc_hd__a21o_1 _4951_ (.A1(_1979_),
    .A2(_2257_),
    .B1(_2266_),
    .X(_0747_));
 sky130_fd_sc_hd__and3_1 _4952_ (.A(_2262_),
    .B(\immu_1.page_table[7][6] ),
    .C(_2259_),
    .X(_2267_));
 sky130_fd_sc_hd__a21o_1 _4953_ (.A1(_1981_),
    .A2(_2257_),
    .B1(_2267_),
    .X(_0748_));
 sky130_fd_sc_hd__and3_1 _4954_ (.A(_2262_),
    .B(\immu_1.page_table[7][7] ),
    .C(_2259_),
    .X(_2268_));
 sky130_fd_sc_hd__a21o_1 _4955_ (.A1(_1983_),
    .A2(_2257_),
    .B1(_2268_),
    .X(_0749_));
 sky130_fd_sc_hd__and3_1 _4956_ (.A(_2262_),
    .B(\immu_1.page_table[7][8] ),
    .C(_2259_),
    .X(_2269_));
 sky130_fd_sc_hd__a21o_1 _4957_ (.A1(_1985_),
    .A2(_2257_),
    .B1(_2269_),
    .X(_0750_));
 sky130_fd_sc_hd__and3_1 _4958_ (.A(_2262_),
    .B(\immu_1.page_table[7][9] ),
    .C(_2259_),
    .X(_2270_));
 sky130_fd_sc_hd__a21o_1 _4959_ (.A1(_1987_),
    .A2(_2257_),
    .B1(_2270_),
    .X(_0751_));
 sky130_fd_sc_hd__and3_1 _4960_ (.A(_2262_),
    .B(\immu_1.page_table[7][10] ),
    .C(_2258_),
    .X(_2271_));
 sky130_fd_sc_hd__a21o_1 _4961_ (.A1(_1989_),
    .A2(_2256_),
    .B1(_2271_),
    .X(_0752_));
 sky130_fd_sc_hd__or4_4 _4962_ (.A(net188),
    .B(net181),
    .C(net190),
    .D(net189),
    .X(_2272_));
 sky130_fd_sc_hd__or2_1 _4963_ (.A(_1999_),
    .B(_2272_),
    .X(_2273_));
 sky130_fd_sc_hd__buf_4 _4964_ (.A(_2273_),
    .X(_2274_));
 sky130_fd_sc_hd__nand2_1 _4965_ (.A(_2190_),
    .B(_2273_),
    .Y(_2275_));
 sky130_fd_sc_hd__clkinv_2 _4966_ (.A(_2275_),
    .Y(_2276_));
 sky130_fd_sc_hd__a2bb2o_1 _4967_ (.A1_N(_1965_),
    .A2_N(_2274_),
    .B1(_2276_),
    .B2(\immu_1.page_table[0][0] ),
    .X(_0753_));
 sky130_fd_sc_hd__buf_4 _4968_ (.A(_2275_),
    .X(_2277_));
 sky130_fd_sc_hd__o22a_1 _4969_ (.A1(_1967_),
    .A2(_2274_),
    .B1(_2277_),
    .B2(\immu_1.page_table[0][1] ),
    .X(_0754_));
 sky130_fd_sc_hd__o22a_1 _4970_ (.A1(_1972_),
    .A2(_2274_),
    .B1(_2277_),
    .B2(\immu_1.page_table[0][2] ),
    .X(_0755_));
 sky130_fd_sc_hd__o22a_1 _4971_ (.A1(_1974_),
    .A2(_2274_),
    .B1(_2277_),
    .B2(\immu_1.page_table[0][3] ),
    .X(_0756_));
 sky130_fd_sc_hd__o22a_1 _4972_ (.A1(_1977_),
    .A2(_2274_),
    .B1(_2277_),
    .B2(\immu_1.page_table[0][4] ),
    .X(_0757_));
 sky130_fd_sc_hd__o22a_1 _4973_ (.A1(_1979_),
    .A2(_2274_),
    .B1(_2277_),
    .B2(\immu_1.page_table[0][5] ),
    .X(_0758_));
 sky130_fd_sc_hd__o22a_1 _4974_ (.A1(_1981_),
    .A2(_2274_),
    .B1(_2277_),
    .B2(\immu_1.page_table[0][6] ),
    .X(_0759_));
 sky130_fd_sc_hd__o22a_1 _4975_ (.A1(_1983_),
    .A2(_2274_),
    .B1(_2277_),
    .B2(\immu_1.page_table[0][7] ),
    .X(_0760_));
 sky130_fd_sc_hd__o22a_1 _4976_ (.A1(_1985_),
    .A2(_2274_),
    .B1(_2277_),
    .B2(\immu_1.page_table[0][8] ),
    .X(_0761_));
 sky130_fd_sc_hd__o22a_1 _4977_ (.A1(_1987_),
    .A2(_2274_),
    .B1(_2277_),
    .B2(\immu_1.page_table[0][9] ),
    .X(_0762_));
 sky130_fd_sc_hd__o22a_1 _4978_ (.A1(_1989_),
    .A2(_2273_),
    .B1(_2277_),
    .B2(\immu_1.page_table[0][10] ),
    .X(_0763_));
 sky130_fd_sc_hd__or2_2 _4979_ (.A(_1960_),
    .B(_2063_),
    .X(_2278_));
 sky130_fd_sc_hd__nor2_1 _4980_ (.A(_1999_),
    .B(_2278_),
    .Y(_2279_));
 sky130_fd_sc_hd__clkbuf_4 _4981_ (.A(_2279_),
    .X(_2280_));
 sky130_fd_sc_hd__or2_1 _4982_ (.A(_2084_),
    .B(_2278_),
    .X(_2281_));
 sky130_fd_sc_hd__buf_2 _4983_ (.A(_2281_),
    .X(_2282_));
 sky130_fd_sc_hd__and3_1 _4984_ (.A(_2262_),
    .B(\immu_1.page_table[15][0] ),
    .C(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__a21o_1 _4985_ (.A1(_1995_),
    .A2(_2280_),
    .B1(_2283_),
    .X(_0764_));
 sky130_fd_sc_hd__buf_2 _4986_ (.A(_2105_),
    .X(_2284_));
 sky130_fd_sc_hd__and3_1 _4987_ (.A(_2284_),
    .B(\immu_1.page_table[15][1] ),
    .C(_2282_),
    .X(_2285_));
 sky130_fd_sc_hd__a21o_1 _4988_ (.A1(_1967_),
    .A2(_2280_),
    .B1(_2285_),
    .X(_0765_));
 sky130_fd_sc_hd__and3_1 _4989_ (.A(_2284_),
    .B(\immu_1.page_table[15][2] ),
    .C(_2282_),
    .X(_2286_));
 sky130_fd_sc_hd__a21o_1 _4990_ (.A1(_1972_),
    .A2(_2280_),
    .B1(_2286_),
    .X(_0766_));
 sky130_fd_sc_hd__and3_1 _4991_ (.A(_2284_),
    .B(\immu_1.page_table[15][3] ),
    .C(_2282_),
    .X(_2287_));
 sky130_fd_sc_hd__a21o_1 _4992_ (.A1(_1974_),
    .A2(_2280_),
    .B1(_2287_),
    .X(_0767_));
 sky130_fd_sc_hd__and3_1 _4993_ (.A(_2284_),
    .B(\immu_1.page_table[15][4] ),
    .C(_2282_),
    .X(_2288_));
 sky130_fd_sc_hd__a21o_1 _4994_ (.A1(_1977_),
    .A2(_2280_),
    .B1(_2288_),
    .X(_0768_));
 sky130_fd_sc_hd__and3_1 _4995_ (.A(_2284_),
    .B(\immu_1.page_table[15][5] ),
    .C(_2282_),
    .X(_2289_));
 sky130_fd_sc_hd__a21o_1 _4996_ (.A1(_1979_),
    .A2(_2280_),
    .B1(_2289_),
    .X(_0769_));
 sky130_fd_sc_hd__and3_1 _4997_ (.A(_2284_),
    .B(\immu_1.page_table[15][6] ),
    .C(_2282_),
    .X(_2290_));
 sky130_fd_sc_hd__a21o_1 _4998_ (.A1(_1981_),
    .A2(_2280_),
    .B1(_2290_),
    .X(_0770_));
 sky130_fd_sc_hd__and3_1 _4999_ (.A(_2284_),
    .B(\immu_1.page_table[15][7] ),
    .C(_2282_),
    .X(_2291_));
 sky130_fd_sc_hd__a21o_1 _5000_ (.A1(_1983_),
    .A2(_2280_),
    .B1(_2291_),
    .X(_0771_));
 sky130_fd_sc_hd__and3_1 _5001_ (.A(_2284_),
    .B(\immu_1.page_table[15][8] ),
    .C(_2282_),
    .X(_2292_));
 sky130_fd_sc_hd__a21o_1 _5002_ (.A1(_1985_),
    .A2(_2280_),
    .B1(_2292_),
    .X(_0772_));
 sky130_fd_sc_hd__and3_1 _5003_ (.A(_2284_),
    .B(\immu_1.page_table[15][9] ),
    .C(_2282_),
    .X(_2293_));
 sky130_fd_sc_hd__a21o_1 _5004_ (.A1(_1987_),
    .A2(_2280_),
    .B1(_2293_),
    .X(_0773_));
 sky130_fd_sc_hd__and3_1 _5005_ (.A(_2284_),
    .B(\immu_1.page_table[15][10] ),
    .C(_2281_),
    .X(_2294_));
 sky130_fd_sc_hd__a21o_1 _5006_ (.A1(_1989_),
    .A2(_2279_),
    .B1(_2294_),
    .X(_0774_));
 sky130_fd_sc_hd__nand2_1 _5007_ (.A(net85),
    .B(net84),
    .Y(_2295_));
 sky130_fd_sc_hd__or2_4 _5008_ (.A(_1912_),
    .B(_2295_),
    .X(_2296_));
 sky130_fd_sc_hd__or2_1 _5009_ (.A(_1922_),
    .B(_2296_),
    .X(_2297_));
 sky130_fd_sc_hd__clkbuf_4 _5010_ (.A(_2297_),
    .X(_2298_));
 sky130_fd_sc_hd__nor2_1 _5011_ (.A(_1926_),
    .B(_2297_),
    .Y(_2299_));
 sky130_fd_sc_hd__a31o_1 _5012_ (.A1(_1976_),
    .A2(\immu_0.page_table[15][0] ),
    .A3(_2298_),
    .B1(_2299_),
    .X(_0775_));
 sky130_fd_sc_hd__buf_4 _5013_ (.A(_1897_),
    .X(_2300_));
 sky130_fd_sc_hd__clkbuf_4 _5014_ (.A(_2300_),
    .X(_2301_));
 sky130_fd_sc_hd__nor2_4 _5015_ (.A(_1930_),
    .B(_2296_),
    .Y(_2302_));
 sky130_fd_sc_hd__and2_1 _5016_ (.A(_1928_),
    .B(_2302_),
    .X(_2303_));
 sky130_fd_sc_hd__a31o_1 _5017_ (.A1(_2301_),
    .A2(\immu_0.page_table[15][1] ),
    .A3(_2298_),
    .B1(_2303_),
    .X(_0776_));
 sky130_fd_sc_hd__and2_1 _5018_ (.A(_1933_),
    .B(_2302_),
    .X(_2304_));
 sky130_fd_sc_hd__a31o_1 _5019_ (.A1(_2301_),
    .A2(\immu_0.page_table[15][2] ),
    .A3(_2298_),
    .B1(_2304_),
    .X(_0777_));
 sky130_fd_sc_hd__and2_1 _5020_ (.A(_1935_),
    .B(_2302_),
    .X(_2305_));
 sky130_fd_sc_hd__a31o_1 _5021_ (.A1(_2301_),
    .A2(\immu_0.page_table[15][3] ),
    .A3(_2298_),
    .B1(_2305_),
    .X(_0778_));
 sky130_fd_sc_hd__and2_1 _5022_ (.A(_1937_),
    .B(_2302_),
    .X(_2306_));
 sky130_fd_sc_hd__a31o_1 _5023_ (.A1(_2301_),
    .A2(\immu_0.page_table[15][4] ),
    .A3(_2298_),
    .B1(_2306_),
    .X(_0779_));
 sky130_fd_sc_hd__and2_1 _5024_ (.A(_1940_),
    .B(_2302_),
    .X(_2307_));
 sky130_fd_sc_hd__a31o_1 _5025_ (.A1(_2301_),
    .A2(\immu_0.page_table[15][5] ),
    .A3(_2298_),
    .B1(_2307_),
    .X(_0780_));
 sky130_fd_sc_hd__and2_1 _5026_ (.A(_1942_),
    .B(_2302_),
    .X(_2308_));
 sky130_fd_sc_hd__a31o_1 _5027_ (.A1(_2301_),
    .A2(\immu_0.page_table[15][6] ),
    .A3(_2298_),
    .B1(_2308_),
    .X(_0781_));
 sky130_fd_sc_hd__and2_1 _5028_ (.A(_1944_),
    .B(_2302_),
    .X(_2309_));
 sky130_fd_sc_hd__a31o_1 _5029_ (.A1(_2301_),
    .A2(\immu_0.page_table[15][7] ),
    .A3(_2298_),
    .B1(_2309_),
    .X(_0782_));
 sky130_fd_sc_hd__buf_4 _5030_ (.A(net103),
    .X(_2310_));
 sky130_fd_sc_hd__and2_1 _5031_ (.A(_2310_),
    .B(_2302_),
    .X(_2311_));
 sky130_fd_sc_hd__a31o_1 _5032_ (.A1(_2301_),
    .A2(\immu_0.page_table[15][8] ),
    .A3(_2298_),
    .B1(_2311_),
    .X(_0783_));
 sky130_fd_sc_hd__buf_4 _5033_ (.A(net104),
    .X(_2312_));
 sky130_fd_sc_hd__and2_1 _5034_ (.A(_2312_),
    .B(_2302_),
    .X(_2313_));
 sky130_fd_sc_hd__a31o_1 _5035_ (.A1(_2301_),
    .A2(\immu_0.page_table[15][9] ),
    .A3(_2298_),
    .B1(_2313_),
    .X(_0784_));
 sky130_fd_sc_hd__buf_4 _5036_ (.A(net93),
    .X(_2314_));
 sky130_fd_sc_hd__and2_1 _5037_ (.A(_2314_),
    .B(_2302_),
    .X(_2315_));
 sky130_fd_sc_hd__a31o_1 _5038_ (.A1(_2301_),
    .A2(\immu_0.page_table[15][10] ),
    .A3(_2297_),
    .B1(_2315_),
    .X(_0785_));
 sky130_fd_sc_hd__clkbuf_4 _5039_ (.A(_2300_),
    .X(_2316_));
 sky130_fd_sc_hd__or2b_1 _5040_ (.A(net76),
    .B_N(net83),
    .X(_2317_));
 sky130_fd_sc_hd__or2_4 _5041_ (.A(_2295_),
    .B(_2317_),
    .X(_2318_));
 sky130_fd_sc_hd__or2_1 _5042_ (.A(_1922_),
    .B(_2318_),
    .X(_2319_));
 sky130_fd_sc_hd__clkbuf_4 _5043_ (.A(_2319_),
    .X(_2320_));
 sky130_fd_sc_hd__nor2_1 _5044_ (.A(_1926_),
    .B(_2319_),
    .Y(_2321_));
 sky130_fd_sc_hd__a31o_1 _5045_ (.A1(_2316_),
    .A2(\immu_0.page_table[14][0] ),
    .A3(_2320_),
    .B1(_2321_),
    .X(_0786_));
 sky130_fd_sc_hd__nor2_4 _5046_ (.A(_1930_),
    .B(_2318_),
    .Y(_2322_));
 sky130_fd_sc_hd__and2_1 _5047_ (.A(_1928_),
    .B(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__a31o_1 _5048_ (.A1(_2316_),
    .A2(\immu_0.page_table[14][1] ),
    .A3(_2320_),
    .B1(_2323_),
    .X(_0787_));
 sky130_fd_sc_hd__and2_1 _5049_ (.A(_1933_),
    .B(_2322_),
    .X(_2324_));
 sky130_fd_sc_hd__a31o_1 _5050_ (.A1(_2316_),
    .A2(\immu_0.page_table[14][2] ),
    .A3(_2320_),
    .B1(_2324_),
    .X(_0788_));
 sky130_fd_sc_hd__and2_1 _5051_ (.A(_1935_),
    .B(_2322_),
    .X(_2325_));
 sky130_fd_sc_hd__a31o_1 _5052_ (.A1(_2316_),
    .A2(\immu_0.page_table[14][3] ),
    .A3(_2320_),
    .B1(_2325_),
    .X(_0789_));
 sky130_fd_sc_hd__and2_1 _5053_ (.A(_1937_),
    .B(_2322_),
    .X(_2326_));
 sky130_fd_sc_hd__a31o_1 _5054_ (.A1(_2316_),
    .A2(\immu_0.page_table[14][4] ),
    .A3(_2320_),
    .B1(_2326_),
    .X(_0790_));
 sky130_fd_sc_hd__and2_1 _5055_ (.A(_1940_),
    .B(_2322_),
    .X(_2327_));
 sky130_fd_sc_hd__a31o_1 _5056_ (.A1(_2316_),
    .A2(\immu_0.page_table[14][5] ),
    .A3(_2320_),
    .B1(_2327_),
    .X(_0791_));
 sky130_fd_sc_hd__and2_1 _5057_ (.A(_1942_),
    .B(_2322_),
    .X(_2328_));
 sky130_fd_sc_hd__a31o_1 _5058_ (.A1(_2316_),
    .A2(\immu_0.page_table[14][6] ),
    .A3(_2320_),
    .B1(_2328_),
    .X(_0792_));
 sky130_fd_sc_hd__and2_1 _5059_ (.A(_1944_),
    .B(_2322_),
    .X(_2329_));
 sky130_fd_sc_hd__a31o_1 _5060_ (.A1(_2316_),
    .A2(\immu_0.page_table[14][7] ),
    .A3(_2320_),
    .B1(_2329_),
    .X(_0793_));
 sky130_fd_sc_hd__and2_1 _5061_ (.A(_2310_),
    .B(_2322_),
    .X(_2330_));
 sky130_fd_sc_hd__a31o_1 _5062_ (.A1(_2316_),
    .A2(\immu_0.page_table[14][8] ),
    .A3(_2320_),
    .B1(_2330_),
    .X(_0794_));
 sky130_fd_sc_hd__and2_1 _5063_ (.A(_2312_),
    .B(_2322_),
    .X(_2331_));
 sky130_fd_sc_hd__a31o_1 _5064_ (.A1(_2316_),
    .A2(\immu_0.page_table[14][9] ),
    .A3(_2320_),
    .B1(_2331_),
    .X(_0795_));
 sky130_fd_sc_hd__buf_4 _5065_ (.A(_2300_),
    .X(_2332_));
 sky130_fd_sc_hd__and2_1 _5066_ (.A(_2314_),
    .B(_2322_),
    .X(_2333_));
 sky130_fd_sc_hd__a31o_1 _5067_ (.A1(_2332_),
    .A2(\immu_0.page_table[14][10] ),
    .A3(_2319_),
    .B1(_2333_),
    .X(_0796_));
 sky130_fd_sc_hd__or3_4 _5068_ (.A(net83),
    .B(net76),
    .C(_2295_),
    .X(_2334_));
 sky130_fd_sc_hd__or2_1 _5069_ (.A(_1922_),
    .B(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__clkbuf_4 _5070_ (.A(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__nor2_1 _5071_ (.A(_1926_),
    .B(_2335_),
    .Y(_2337_));
 sky130_fd_sc_hd__a31o_1 _5072_ (.A1(_2332_),
    .A2(\immu_0.page_table[12][0] ),
    .A3(_2336_),
    .B1(_2337_),
    .X(_0797_));
 sky130_fd_sc_hd__nor2_4 _5073_ (.A(_1930_),
    .B(_2334_),
    .Y(_2338_));
 sky130_fd_sc_hd__and2_1 _5074_ (.A(_1928_),
    .B(_2338_),
    .X(_2339_));
 sky130_fd_sc_hd__a31o_1 _5075_ (.A1(_2332_),
    .A2(\immu_0.page_table[12][1] ),
    .A3(_2336_),
    .B1(_2339_),
    .X(_0798_));
 sky130_fd_sc_hd__and2_1 _5076_ (.A(_1933_),
    .B(_2338_),
    .X(_2340_));
 sky130_fd_sc_hd__a31o_1 _5077_ (.A1(_2332_),
    .A2(\immu_0.page_table[12][2] ),
    .A3(_2336_),
    .B1(_2340_),
    .X(_0799_));
 sky130_fd_sc_hd__and2_1 _5078_ (.A(_1935_),
    .B(_2338_),
    .X(_2341_));
 sky130_fd_sc_hd__a31o_1 _5079_ (.A1(_2332_),
    .A2(\immu_0.page_table[12][3] ),
    .A3(_2336_),
    .B1(_2341_),
    .X(_0800_));
 sky130_fd_sc_hd__and2_1 _5080_ (.A(_1937_),
    .B(_2338_),
    .X(_2342_));
 sky130_fd_sc_hd__a31o_1 _5081_ (.A1(_2332_),
    .A2(\immu_0.page_table[12][4] ),
    .A3(_2336_),
    .B1(_2342_),
    .X(_0801_));
 sky130_fd_sc_hd__and2_1 _5082_ (.A(_1940_),
    .B(_2338_),
    .X(_2343_));
 sky130_fd_sc_hd__a31o_1 _5083_ (.A1(_2332_),
    .A2(\immu_0.page_table[12][5] ),
    .A3(_2336_),
    .B1(_2343_),
    .X(_0802_));
 sky130_fd_sc_hd__and2_1 _5084_ (.A(_1942_),
    .B(_2338_),
    .X(_2344_));
 sky130_fd_sc_hd__a31o_1 _5085_ (.A1(_2332_),
    .A2(\immu_0.page_table[12][6] ),
    .A3(_2336_),
    .B1(_2344_),
    .X(_0803_));
 sky130_fd_sc_hd__and2_1 _5086_ (.A(_1944_),
    .B(_2338_),
    .X(_2345_));
 sky130_fd_sc_hd__a31o_1 _5087_ (.A1(_2332_),
    .A2(\immu_0.page_table[12][7] ),
    .A3(_2336_),
    .B1(_2345_),
    .X(_0804_));
 sky130_fd_sc_hd__and2_1 _5088_ (.A(_2310_),
    .B(_2338_),
    .X(_2346_));
 sky130_fd_sc_hd__a31o_1 _5089_ (.A1(_2332_),
    .A2(\immu_0.page_table[12][8] ),
    .A3(_2336_),
    .B1(_2346_),
    .X(_0805_));
 sky130_fd_sc_hd__clkbuf_4 _5090_ (.A(_2300_),
    .X(_2347_));
 sky130_fd_sc_hd__and2_1 _5091_ (.A(_2312_),
    .B(_2338_),
    .X(_2348_));
 sky130_fd_sc_hd__a31o_1 _5092_ (.A1(_2347_),
    .A2(\immu_0.page_table[12][9] ),
    .A3(_2336_),
    .B1(_2348_),
    .X(_0806_));
 sky130_fd_sc_hd__and2_1 _5093_ (.A(_2314_),
    .B(_2338_),
    .X(_2349_));
 sky130_fd_sc_hd__a31o_1 _5094_ (.A1(_2347_),
    .A2(\immu_0.page_table[12][10] ),
    .A3(_2335_),
    .B1(_2349_),
    .X(_0807_));
 sky130_fd_sc_hd__or2b_2 _5095_ (.A(net83),
    .B_N(net76),
    .X(_2350_));
 sky130_fd_sc_hd__or2_4 _5096_ (.A(_2295_),
    .B(_2350_),
    .X(_2351_));
 sky130_fd_sc_hd__or2_1 _5097_ (.A(_1922_),
    .B(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__clkbuf_4 _5098_ (.A(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__nor2_1 _5099_ (.A(_1926_),
    .B(_2352_),
    .Y(_2354_));
 sky130_fd_sc_hd__a31o_1 _5100_ (.A1(_2347_),
    .A2(\immu_0.page_table[13][0] ),
    .A3(_2353_),
    .B1(_2354_),
    .X(_0808_));
 sky130_fd_sc_hd__nor2_4 _5101_ (.A(_1930_),
    .B(_2351_),
    .Y(_2355_));
 sky130_fd_sc_hd__and2_1 _5102_ (.A(_1928_),
    .B(_2355_),
    .X(_2356_));
 sky130_fd_sc_hd__a31o_1 _5103_ (.A1(_2347_),
    .A2(\immu_0.page_table[13][1] ),
    .A3(_2353_),
    .B1(_2356_),
    .X(_0000_));
 sky130_fd_sc_hd__and2_1 _5104_ (.A(_1933_),
    .B(_2355_),
    .X(_2357_));
 sky130_fd_sc_hd__a31o_1 _5105_ (.A1(_2347_),
    .A2(\immu_0.page_table[13][2] ),
    .A3(_2353_),
    .B1(_2357_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _5106_ (.A(_1935_),
    .B(_2355_),
    .X(_2358_));
 sky130_fd_sc_hd__a31o_1 _5107_ (.A1(_2347_),
    .A2(\immu_0.page_table[13][3] ),
    .A3(_2353_),
    .B1(_2358_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _5108_ (.A(_1937_),
    .B(_2355_),
    .X(_2359_));
 sky130_fd_sc_hd__a31o_1 _5109_ (.A1(_2347_),
    .A2(\immu_0.page_table[13][4] ),
    .A3(_2353_),
    .B1(_2359_),
    .X(_0003_));
 sky130_fd_sc_hd__and2_1 _5110_ (.A(_1940_),
    .B(_2355_),
    .X(_2360_));
 sky130_fd_sc_hd__a31o_1 _5111_ (.A1(_2347_),
    .A2(\immu_0.page_table[13][5] ),
    .A3(_2353_),
    .B1(_2360_),
    .X(_0004_));
 sky130_fd_sc_hd__and2_1 _5112_ (.A(_1942_),
    .B(_2355_),
    .X(_2361_));
 sky130_fd_sc_hd__a31o_1 _5113_ (.A1(_2347_),
    .A2(\immu_0.page_table[13][6] ),
    .A3(_2353_),
    .B1(_2361_),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _5114_ (.A(_1944_),
    .B(_2355_),
    .X(_2362_));
 sky130_fd_sc_hd__a31o_1 _5115_ (.A1(_2347_),
    .A2(\immu_0.page_table[13][7] ),
    .A3(_2353_),
    .B1(_2362_),
    .X(_0006_));
 sky130_fd_sc_hd__buf_4 _5116_ (.A(_2300_),
    .X(_2363_));
 sky130_fd_sc_hd__and2_1 _5117_ (.A(_2310_),
    .B(_2355_),
    .X(_2364_));
 sky130_fd_sc_hd__a31o_1 _5118_ (.A1(_2363_),
    .A2(\immu_0.page_table[13][8] ),
    .A3(_2353_),
    .B1(_2364_),
    .X(_0007_));
 sky130_fd_sc_hd__and2_1 _5119_ (.A(_2312_),
    .B(_2355_),
    .X(_2365_));
 sky130_fd_sc_hd__a31o_1 _5120_ (.A1(_2363_),
    .A2(\immu_0.page_table[13][9] ),
    .A3(_2353_),
    .B1(_2365_),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _5121_ (.A(_2314_),
    .B(_2355_),
    .X(_2366_));
 sky130_fd_sc_hd__a31o_1 _5122_ (.A1(_2363_),
    .A2(\immu_0.page_table[13][10] ),
    .A3(_2352_),
    .B1(_2366_),
    .X(_0009_));
 sky130_fd_sc_hd__or2_4 _5123_ (.A(_1913_),
    .B(_2317_),
    .X(_2367_));
 sky130_fd_sc_hd__nor2_1 _5124_ (.A(_2217_),
    .B(_2367_),
    .Y(_2368_));
 sky130_fd_sc_hd__buf_4 _5125_ (.A(_2368_),
    .X(_2369_));
 sky130_fd_sc_hd__buf_2 _5126_ (.A(_1896_),
    .X(_2370_));
 sky130_fd_sc_hd__buf_2 _5127_ (.A(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__or2_1 _5128_ (.A(_2216_),
    .B(_2367_),
    .X(_2372_));
 sky130_fd_sc_hd__clkbuf_4 _5129_ (.A(_2372_),
    .X(_2373_));
 sky130_fd_sc_hd__and3_1 _5130_ (.A(_2371_),
    .B(\dmmu0.page_table[10][0] ),
    .C(_2373_),
    .X(_2374_));
 sky130_fd_sc_hd__a21o_1 _5131_ (.A1(_2211_),
    .A2(_2369_),
    .B1(_2374_),
    .X(_0010_));
 sky130_fd_sc_hd__and3_1 _5132_ (.A(_2371_),
    .B(\dmmu0.page_table[10][1] ),
    .C(_2373_),
    .X(_2375_));
 sky130_fd_sc_hd__a21o_1 _5133_ (.A1(_2224_),
    .A2(_2369_),
    .B1(_2375_),
    .X(_0011_));
 sky130_fd_sc_hd__and3_1 _5134_ (.A(_2371_),
    .B(\dmmu0.page_table[10][2] ),
    .C(_2373_),
    .X(_2376_));
 sky130_fd_sc_hd__a21o_1 _5135_ (.A1(_2227_),
    .A2(_2369_),
    .B1(_2376_),
    .X(_0012_));
 sky130_fd_sc_hd__and3_1 _5136_ (.A(_2371_),
    .B(\dmmu0.page_table[10][3] ),
    .C(_2373_),
    .X(_2377_));
 sky130_fd_sc_hd__a21o_1 _5137_ (.A1(_2230_),
    .A2(_2369_),
    .B1(_2377_),
    .X(_0013_));
 sky130_fd_sc_hd__and3_1 _5138_ (.A(_2371_),
    .B(\dmmu0.page_table[10][4] ),
    .C(_2373_),
    .X(_2378_));
 sky130_fd_sc_hd__a21o_1 _5139_ (.A1(_2233_),
    .A2(_2369_),
    .B1(_2378_),
    .X(_0014_));
 sky130_fd_sc_hd__and3_1 _5140_ (.A(_2371_),
    .B(\dmmu0.page_table[10][5] ),
    .C(_2373_),
    .X(_2379_));
 sky130_fd_sc_hd__a21o_1 _5141_ (.A1(_2236_),
    .A2(_2369_),
    .B1(_2379_),
    .X(_0015_));
 sky130_fd_sc_hd__and3_1 _5142_ (.A(_2371_),
    .B(\dmmu0.page_table[10][6] ),
    .C(_2373_),
    .X(_2380_));
 sky130_fd_sc_hd__a21o_1 _5143_ (.A1(_2240_),
    .A2(_2369_),
    .B1(_2380_),
    .X(_0016_));
 sky130_fd_sc_hd__and3_1 _5144_ (.A(_2371_),
    .B(\dmmu0.page_table[10][7] ),
    .C(_2373_),
    .X(_2381_));
 sky130_fd_sc_hd__a21o_1 _5145_ (.A1(_2243_),
    .A2(_2369_),
    .B1(_2381_),
    .X(_0017_));
 sky130_fd_sc_hd__and3_1 _5146_ (.A(_2371_),
    .B(\dmmu0.page_table[10][8] ),
    .C(_2373_),
    .X(_2382_));
 sky130_fd_sc_hd__a21o_1 _5147_ (.A1(_2245_),
    .A2(_2369_),
    .B1(_2382_),
    .X(_0018_));
 sky130_fd_sc_hd__and3_1 _5148_ (.A(_2371_),
    .B(\dmmu0.page_table[10][9] ),
    .C(_2373_),
    .X(_2383_));
 sky130_fd_sc_hd__a21o_1 _5149_ (.A1(_2247_),
    .A2(_2369_),
    .B1(_2383_),
    .X(_0019_));
 sky130_fd_sc_hd__buf_2 _5150_ (.A(_2370_),
    .X(_2384_));
 sky130_fd_sc_hd__and3_1 _5151_ (.A(_2384_),
    .B(\dmmu0.page_table[10][10] ),
    .C(_2372_),
    .X(_2385_));
 sky130_fd_sc_hd__a21o_1 _5152_ (.A1(_2249_),
    .A2(_2368_),
    .B1(_2385_),
    .X(_0020_));
 sky130_fd_sc_hd__and3_1 _5153_ (.A(_2384_),
    .B(\dmmu0.page_table[10][11] ),
    .C(_2372_),
    .X(_2386_));
 sky130_fd_sc_hd__a21o_1 _5154_ (.A1(_2251_),
    .A2(_2368_),
    .B1(_2386_),
    .X(_0021_));
 sky130_fd_sc_hd__and3_1 _5155_ (.A(_2384_),
    .B(\dmmu0.page_table[10][12] ),
    .C(_2372_),
    .X(_2387_));
 sky130_fd_sc_hd__a21o_1 _5156_ (.A1(_2253_),
    .A2(_2368_),
    .B1(_2387_),
    .X(_0022_));
 sky130_fd_sc_hd__or2_4 _5157_ (.A(_1913_),
    .B(_2350_),
    .X(_2388_));
 sky130_fd_sc_hd__nor2_1 _5158_ (.A(_2217_),
    .B(_2388_),
    .Y(_2389_));
 sky130_fd_sc_hd__buf_4 _5159_ (.A(_2389_),
    .X(_2390_));
 sky130_fd_sc_hd__or2_1 _5160_ (.A(_2216_),
    .B(_2388_),
    .X(_2391_));
 sky130_fd_sc_hd__clkbuf_4 _5161_ (.A(_2391_),
    .X(_2392_));
 sky130_fd_sc_hd__and3_1 _5162_ (.A(_2384_),
    .B(\dmmu0.page_table[9][0] ),
    .C(_2392_),
    .X(_2393_));
 sky130_fd_sc_hd__a21o_1 _5163_ (.A1(_2211_),
    .A2(_2390_),
    .B1(_2393_),
    .X(_0023_));
 sky130_fd_sc_hd__and3_1 _5164_ (.A(_2384_),
    .B(\dmmu0.page_table[9][1] ),
    .C(_2392_),
    .X(_2394_));
 sky130_fd_sc_hd__a21o_1 _5165_ (.A1(_2224_),
    .A2(_2390_),
    .B1(_2394_),
    .X(_0024_));
 sky130_fd_sc_hd__and3_1 _5166_ (.A(_2384_),
    .B(\dmmu0.page_table[9][2] ),
    .C(_2392_),
    .X(_2395_));
 sky130_fd_sc_hd__a21o_1 _5167_ (.A1(_2227_),
    .A2(_2390_),
    .B1(_2395_),
    .X(_0025_));
 sky130_fd_sc_hd__and3_1 _5168_ (.A(_2384_),
    .B(\dmmu0.page_table[9][3] ),
    .C(_2392_),
    .X(_2396_));
 sky130_fd_sc_hd__a21o_1 _5169_ (.A1(_2230_),
    .A2(_2390_),
    .B1(_2396_),
    .X(_0026_));
 sky130_fd_sc_hd__and3_1 _5170_ (.A(_2384_),
    .B(\dmmu0.page_table[9][4] ),
    .C(_2392_),
    .X(_2397_));
 sky130_fd_sc_hd__a21o_1 _5171_ (.A1(_2233_),
    .A2(_2390_),
    .B1(_2397_),
    .X(_0027_));
 sky130_fd_sc_hd__and3_1 _5172_ (.A(_2384_),
    .B(\dmmu0.page_table[9][5] ),
    .C(_2392_),
    .X(_2398_));
 sky130_fd_sc_hd__a21o_1 _5173_ (.A1(_2236_),
    .A2(_2390_),
    .B1(_2398_),
    .X(_0028_));
 sky130_fd_sc_hd__and3_1 _5174_ (.A(_2384_),
    .B(\dmmu0.page_table[9][6] ),
    .C(_2392_),
    .X(_2399_));
 sky130_fd_sc_hd__a21o_1 _5175_ (.A1(_2240_),
    .A2(_2390_),
    .B1(_2399_),
    .X(_0029_));
 sky130_fd_sc_hd__clkbuf_4 _5176_ (.A(_2370_),
    .X(_2400_));
 sky130_fd_sc_hd__and3_1 _5177_ (.A(_2400_),
    .B(\dmmu0.page_table[9][7] ),
    .C(_2392_),
    .X(_2401_));
 sky130_fd_sc_hd__a21o_1 _5178_ (.A1(_2243_),
    .A2(_2390_),
    .B1(_2401_),
    .X(_0030_));
 sky130_fd_sc_hd__and3_1 _5179_ (.A(_2400_),
    .B(\dmmu0.page_table[9][8] ),
    .C(_2392_),
    .X(_2402_));
 sky130_fd_sc_hd__a21o_1 _5180_ (.A1(_2245_),
    .A2(_2390_),
    .B1(_2402_),
    .X(_0031_));
 sky130_fd_sc_hd__and3_1 _5181_ (.A(_2400_),
    .B(\dmmu0.page_table[9][9] ),
    .C(_2392_),
    .X(_2403_));
 sky130_fd_sc_hd__a21o_1 _5182_ (.A1(_2247_),
    .A2(_2390_),
    .B1(_2403_),
    .X(_0032_));
 sky130_fd_sc_hd__and3_1 _5183_ (.A(_2400_),
    .B(\dmmu0.page_table[9][10] ),
    .C(_2391_),
    .X(_2404_));
 sky130_fd_sc_hd__a21o_1 _5184_ (.A1(_2249_),
    .A2(_2389_),
    .B1(_2404_),
    .X(_0033_));
 sky130_fd_sc_hd__and3_1 _5185_ (.A(_2400_),
    .B(\dmmu0.page_table[9][11] ),
    .C(_2391_),
    .X(_2405_));
 sky130_fd_sc_hd__a21o_1 _5186_ (.A1(_2251_),
    .A2(_2389_),
    .B1(_2405_),
    .X(_0034_));
 sky130_fd_sc_hd__and3_1 _5187_ (.A(_2400_),
    .B(\dmmu0.page_table[9][12] ),
    .C(_2391_),
    .X(_2406_));
 sky130_fd_sc_hd__a21o_1 _5188_ (.A1(_2253_),
    .A2(_2389_),
    .B1(_2406_),
    .X(_0035_));
 sky130_fd_sc_hd__or3_4 _5189_ (.A(net83),
    .B(net76),
    .C(_1913_),
    .X(_2407_));
 sky130_fd_sc_hd__nor2_1 _5190_ (.A(_2217_),
    .B(_2407_),
    .Y(_2408_));
 sky130_fd_sc_hd__buf_4 _5191_ (.A(_2408_),
    .X(_2409_));
 sky130_fd_sc_hd__or2_1 _5192_ (.A(_2216_),
    .B(_2407_),
    .X(_2410_));
 sky130_fd_sc_hd__clkbuf_4 _5193_ (.A(_2410_),
    .X(_2411_));
 sky130_fd_sc_hd__and3_1 _5194_ (.A(_2400_),
    .B(\dmmu0.page_table[8][0] ),
    .C(_2411_),
    .X(_2412_));
 sky130_fd_sc_hd__a21o_1 _5195_ (.A1(_2211_),
    .A2(_2409_),
    .B1(_2412_),
    .X(_0036_));
 sky130_fd_sc_hd__and3_1 _5196_ (.A(_2400_),
    .B(\dmmu0.page_table[8][1] ),
    .C(_2411_),
    .X(_2413_));
 sky130_fd_sc_hd__a21o_1 _5197_ (.A1(_2224_),
    .A2(_2409_),
    .B1(_2413_),
    .X(_0037_));
 sky130_fd_sc_hd__and3_1 _5198_ (.A(_2400_),
    .B(\dmmu0.page_table[8][2] ),
    .C(_2411_),
    .X(_2414_));
 sky130_fd_sc_hd__a21o_1 _5199_ (.A1(_2227_),
    .A2(_2409_),
    .B1(_2414_),
    .X(_0038_));
 sky130_fd_sc_hd__and3_1 _5200_ (.A(_2400_),
    .B(\dmmu0.page_table[8][3] ),
    .C(_2411_),
    .X(_2415_));
 sky130_fd_sc_hd__a21o_1 _5201_ (.A1(_2230_),
    .A2(_2409_),
    .B1(_2415_),
    .X(_0039_));
 sky130_fd_sc_hd__clkbuf_4 _5202_ (.A(_2370_),
    .X(_2416_));
 sky130_fd_sc_hd__and3_1 _5203_ (.A(_2416_),
    .B(\dmmu0.page_table[8][4] ),
    .C(_2411_),
    .X(_2417_));
 sky130_fd_sc_hd__a21o_1 _5204_ (.A1(_2233_),
    .A2(_2409_),
    .B1(_2417_),
    .X(_0040_));
 sky130_fd_sc_hd__and3_1 _5205_ (.A(_2416_),
    .B(\dmmu0.page_table[8][5] ),
    .C(_2411_),
    .X(_2418_));
 sky130_fd_sc_hd__a21o_1 _5206_ (.A1(_2236_),
    .A2(_2409_),
    .B1(_2418_),
    .X(_0041_));
 sky130_fd_sc_hd__and3_1 _5207_ (.A(_2416_),
    .B(\dmmu0.page_table[8][6] ),
    .C(_2411_),
    .X(_2419_));
 sky130_fd_sc_hd__a21o_1 _5208_ (.A1(_2240_),
    .A2(_2409_),
    .B1(_2419_),
    .X(_0042_));
 sky130_fd_sc_hd__and3_1 _5209_ (.A(_2416_),
    .B(\dmmu0.page_table[8][7] ),
    .C(_2411_),
    .X(_2420_));
 sky130_fd_sc_hd__a21o_1 _5210_ (.A1(_2243_),
    .A2(_2409_),
    .B1(_2420_),
    .X(_0043_));
 sky130_fd_sc_hd__and3_1 _5211_ (.A(_2416_),
    .B(\dmmu0.page_table[8][8] ),
    .C(_2411_),
    .X(_2421_));
 sky130_fd_sc_hd__a21o_1 _5212_ (.A1(_2245_),
    .A2(_2409_),
    .B1(_2421_),
    .X(_0044_));
 sky130_fd_sc_hd__and3_1 _5213_ (.A(_2416_),
    .B(\dmmu0.page_table[8][9] ),
    .C(_2411_),
    .X(_2422_));
 sky130_fd_sc_hd__a21o_1 _5214_ (.A1(_2247_),
    .A2(_2409_),
    .B1(_2422_),
    .X(_0045_));
 sky130_fd_sc_hd__and3_1 _5215_ (.A(_2416_),
    .B(\dmmu0.page_table[8][10] ),
    .C(_2410_),
    .X(_2423_));
 sky130_fd_sc_hd__a21o_1 _5216_ (.A1(_2249_),
    .A2(_2408_),
    .B1(_2423_),
    .X(_0046_));
 sky130_fd_sc_hd__and3_1 _5217_ (.A(_2416_),
    .B(\dmmu0.page_table[8][11] ),
    .C(_2410_),
    .X(_2424_));
 sky130_fd_sc_hd__a21o_1 _5218_ (.A1(_2251_),
    .A2(_2408_),
    .B1(_2424_),
    .X(_0047_));
 sky130_fd_sc_hd__and3_1 _5219_ (.A(_2416_),
    .B(\dmmu0.page_table[8][12] ),
    .C(_2410_),
    .X(_2425_));
 sky130_fd_sc_hd__a21o_1 _5220_ (.A1(_2253_),
    .A2(_2408_),
    .B1(_2425_),
    .X(_0048_));
 sky130_fd_sc_hd__or4_1 _5221_ (.A(net78),
    .B(net77),
    .C(net91),
    .D(_2213_),
    .X(_2426_));
 sky130_fd_sc_hd__nor2_1 _5222_ (.A(_1919_),
    .B(_2426_),
    .Y(_2427_));
 sky130_fd_sc_hd__and2b_1 _5223_ (.A_N(_2367_),
    .B(_2427_),
    .X(_2428_));
 sky130_fd_sc_hd__or4_2 _5224_ (.A(net196),
    .B(net195),
    .C(_1953_),
    .D(_1956_),
    .X(_2429_));
 sky130_fd_sc_hd__nor2_2 _5225_ (.A(_2081_),
    .B(_2429_),
    .Y(_2430_));
 sky130_fd_sc_hd__a21bo_1 _5226_ (.A1(net197),
    .A2(_2430_),
    .B1_N(net407),
    .X(_2431_));
 sky130_fd_sc_hd__a21oi_1 _5227_ (.A1(_2210_),
    .A2(_2428_),
    .B1(_2431_),
    .Y(_2432_));
 sky130_fd_sc_hd__nor2_2 _5228_ (.A(_1913_),
    .B(_2350_),
    .Y(_2433_));
 sky130_fd_sc_hd__nor2_2 _5229_ (.A(_2099_),
    .B(_2429_),
    .Y(_2434_));
 sky130_fd_sc_hd__a32o_1 _5230_ (.A1(net92),
    .A2(_2433_),
    .A3(_2427_),
    .B1(_2434_),
    .B2(net197),
    .X(_2435_));
 sky130_fd_sc_hd__o21a_1 _5231_ (.A1(_2432_),
    .A2(_2435_),
    .B1(_1911_),
    .X(_0049_));
 sky130_fd_sc_hd__a21bo_1 _5232_ (.A1(net201),
    .A2(_2430_),
    .B1_N(net408),
    .X(_2436_));
 sky130_fd_sc_hd__a21oi_1 _5233_ (.A1(_2223_),
    .A2(_2428_),
    .B1(_2436_),
    .Y(_2437_));
 sky130_fd_sc_hd__a32o_1 _5234_ (.A1(net96),
    .A2(_2433_),
    .A3(_2427_),
    .B1(_2434_),
    .B2(net201),
    .X(_2438_));
 sky130_fd_sc_hd__o21a_1 _5235_ (.A1(_2437_),
    .A2(_2438_),
    .B1(_1911_),
    .X(_0050_));
 sky130_fd_sc_hd__or2b_1 _5236_ (.A(net85),
    .B_N(net84),
    .X(_2439_));
 sky130_fd_sc_hd__or2_4 _5237_ (.A(_1912_),
    .B(_2439_),
    .X(_2440_));
 sky130_fd_sc_hd__nor2_1 _5238_ (.A(_2217_),
    .B(_2440_),
    .Y(_2441_));
 sky130_fd_sc_hd__clkbuf_4 _5239_ (.A(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__clkbuf_4 _5240_ (.A(_2215_),
    .X(_2443_));
 sky130_fd_sc_hd__or2_1 _5241_ (.A(_2443_),
    .B(_2440_),
    .X(_2444_));
 sky130_fd_sc_hd__clkbuf_4 _5242_ (.A(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__and3_1 _5243_ (.A(_2416_),
    .B(\dmmu0.page_table[7][0] ),
    .C(_2445_),
    .X(_2446_));
 sky130_fd_sc_hd__a21o_1 _5244_ (.A1(_2211_),
    .A2(_2442_),
    .B1(_2446_),
    .X(_0051_));
 sky130_fd_sc_hd__clkbuf_4 _5245_ (.A(_2370_),
    .X(_2447_));
 sky130_fd_sc_hd__and3_1 _5246_ (.A(_2447_),
    .B(\dmmu0.page_table[7][1] ),
    .C(_2445_),
    .X(_2448_));
 sky130_fd_sc_hd__a21o_1 _5247_ (.A1(_2224_),
    .A2(_2442_),
    .B1(_2448_),
    .X(_0052_));
 sky130_fd_sc_hd__and3_1 _5248_ (.A(_2447_),
    .B(\dmmu0.page_table[7][2] ),
    .C(_2445_),
    .X(_2449_));
 sky130_fd_sc_hd__a21o_1 _5249_ (.A1(_2227_),
    .A2(_2442_),
    .B1(_2449_),
    .X(_0053_));
 sky130_fd_sc_hd__and3_1 _5250_ (.A(_2447_),
    .B(\dmmu0.page_table[7][3] ),
    .C(_2445_),
    .X(_2450_));
 sky130_fd_sc_hd__a21o_1 _5251_ (.A1(_2230_),
    .A2(_2442_),
    .B1(_2450_),
    .X(_0054_));
 sky130_fd_sc_hd__and3_1 _5252_ (.A(_2447_),
    .B(\dmmu0.page_table[7][4] ),
    .C(_2445_),
    .X(_2451_));
 sky130_fd_sc_hd__a21o_1 _5253_ (.A1(_2233_),
    .A2(_2442_),
    .B1(_2451_),
    .X(_0055_));
 sky130_fd_sc_hd__and3_1 _5254_ (.A(_2447_),
    .B(\dmmu0.page_table[7][5] ),
    .C(_2445_),
    .X(_2452_));
 sky130_fd_sc_hd__a21o_1 _5255_ (.A1(_2236_),
    .A2(_2442_),
    .B1(_2452_),
    .X(_0056_));
 sky130_fd_sc_hd__and3_1 _5256_ (.A(_2447_),
    .B(\dmmu0.page_table[7][6] ),
    .C(_2445_),
    .X(_2453_));
 sky130_fd_sc_hd__a21o_1 _5257_ (.A1(_2240_),
    .A2(_2442_),
    .B1(_2453_),
    .X(_0057_));
 sky130_fd_sc_hd__and3_1 _5258_ (.A(_2447_),
    .B(\dmmu0.page_table[7][7] ),
    .C(_2445_),
    .X(_2454_));
 sky130_fd_sc_hd__a21o_1 _5259_ (.A1(_2243_),
    .A2(_2442_),
    .B1(_2454_),
    .X(_0058_));
 sky130_fd_sc_hd__and3_1 _5260_ (.A(_2447_),
    .B(\dmmu0.page_table[7][8] ),
    .C(_2445_),
    .X(_2455_));
 sky130_fd_sc_hd__a21o_1 _5261_ (.A1(_2245_),
    .A2(_2442_),
    .B1(_2455_),
    .X(_0059_));
 sky130_fd_sc_hd__and3_1 _5262_ (.A(_2447_),
    .B(\dmmu0.page_table[7][9] ),
    .C(_2445_),
    .X(_2456_));
 sky130_fd_sc_hd__a21o_1 _5263_ (.A1(_2247_),
    .A2(_2442_),
    .B1(_2456_),
    .X(_0060_));
 sky130_fd_sc_hd__and3_1 _5264_ (.A(_2447_),
    .B(\dmmu0.page_table[7][10] ),
    .C(_2444_),
    .X(_2457_));
 sky130_fd_sc_hd__a21o_1 _5265_ (.A1(_2249_),
    .A2(_2441_),
    .B1(_2457_),
    .X(_0061_));
 sky130_fd_sc_hd__clkbuf_4 _5266_ (.A(_2370_),
    .X(_2458_));
 sky130_fd_sc_hd__and3_1 _5267_ (.A(_2458_),
    .B(\dmmu0.page_table[7][11] ),
    .C(_2444_),
    .X(_2459_));
 sky130_fd_sc_hd__a21o_1 _5268_ (.A1(_2251_),
    .A2(_2441_),
    .B1(_2459_),
    .X(_0062_));
 sky130_fd_sc_hd__and3_1 _5269_ (.A(_2458_),
    .B(\dmmu0.page_table[7][12] ),
    .C(_2444_),
    .X(_2460_));
 sky130_fd_sc_hd__a21o_1 _5270_ (.A1(_2253_),
    .A2(_2441_),
    .B1(_2460_),
    .X(_0063_));
 sky130_fd_sc_hd__nor2_1 _5271_ (.A(_2217_),
    .B(_2318_),
    .Y(_2461_));
 sky130_fd_sc_hd__buf_4 _5272_ (.A(_2461_),
    .X(_2462_));
 sky130_fd_sc_hd__or2_1 _5273_ (.A(_2443_),
    .B(_2318_),
    .X(_2463_));
 sky130_fd_sc_hd__clkbuf_4 _5274_ (.A(_2463_),
    .X(_2464_));
 sky130_fd_sc_hd__and3_1 _5275_ (.A(_2458_),
    .B(\dmmu0.page_table[14][0] ),
    .C(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__a21o_1 _5276_ (.A1(_2211_),
    .A2(_2462_),
    .B1(_2465_),
    .X(_0064_));
 sky130_fd_sc_hd__and3_1 _5277_ (.A(_2458_),
    .B(\dmmu0.page_table[14][1] ),
    .C(_2464_),
    .X(_2466_));
 sky130_fd_sc_hd__a21o_1 _5278_ (.A1(_2224_),
    .A2(_2462_),
    .B1(_2466_),
    .X(_0065_));
 sky130_fd_sc_hd__and3_1 _5279_ (.A(_2458_),
    .B(\dmmu0.page_table[14][2] ),
    .C(_2464_),
    .X(_2467_));
 sky130_fd_sc_hd__a21o_1 _5280_ (.A1(_2227_),
    .A2(_2462_),
    .B1(_2467_),
    .X(_0066_));
 sky130_fd_sc_hd__and3_1 _5281_ (.A(_2458_),
    .B(\dmmu0.page_table[14][3] ),
    .C(_2464_),
    .X(_2468_));
 sky130_fd_sc_hd__a21o_1 _5282_ (.A1(_2230_),
    .A2(_2462_),
    .B1(_2468_),
    .X(_0067_));
 sky130_fd_sc_hd__and3_1 _5283_ (.A(_2458_),
    .B(\dmmu0.page_table[14][4] ),
    .C(_2464_),
    .X(_2469_));
 sky130_fd_sc_hd__a21o_1 _5284_ (.A1(_2233_),
    .A2(_2462_),
    .B1(_2469_),
    .X(_0068_));
 sky130_fd_sc_hd__and3_1 _5285_ (.A(_2458_),
    .B(\dmmu0.page_table[14][5] ),
    .C(_2464_),
    .X(_2470_));
 sky130_fd_sc_hd__a21o_1 _5286_ (.A1(_2236_),
    .A2(_2462_),
    .B1(_2470_),
    .X(_0069_));
 sky130_fd_sc_hd__and3_1 _5287_ (.A(_2458_),
    .B(\dmmu0.page_table[14][6] ),
    .C(_2464_),
    .X(_2471_));
 sky130_fd_sc_hd__a21o_1 _5288_ (.A1(_2240_),
    .A2(_2462_),
    .B1(_2471_),
    .X(_0070_));
 sky130_fd_sc_hd__and3_1 _5289_ (.A(_2458_),
    .B(\dmmu0.page_table[14][7] ),
    .C(_2464_),
    .X(_2472_));
 sky130_fd_sc_hd__a21o_1 _5290_ (.A1(_2243_),
    .A2(_2462_),
    .B1(_2472_),
    .X(_0071_));
 sky130_fd_sc_hd__clkbuf_4 _5291_ (.A(_2370_),
    .X(_2473_));
 sky130_fd_sc_hd__and3_1 _5292_ (.A(_2473_),
    .B(\dmmu0.page_table[14][8] ),
    .C(_2464_),
    .X(_2474_));
 sky130_fd_sc_hd__a21o_1 _5293_ (.A1(_2245_),
    .A2(_2462_),
    .B1(_2474_),
    .X(_0072_));
 sky130_fd_sc_hd__and3_1 _5294_ (.A(_2473_),
    .B(\dmmu0.page_table[14][9] ),
    .C(_2464_),
    .X(_2475_));
 sky130_fd_sc_hd__a21o_1 _5295_ (.A1(_2247_),
    .A2(_2462_),
    .B1(_2475_),
    .X(_0073_));
 sky130_fd_sc_hd__and3_1 _5296_ (.A(_2473_),
    .B(\dmmu0.page_table[14][10] ),
    .C(_2463_),
    .X(_2476_));
 sky130_fd_sc_hd__a21o_1 _5297_ (.A1(_2249_),
    .A2(_2461_),
    .B1(_2476_),
    .X(_0074_));
 sky130_fd_sc_hd__and3_1 _5298_ (.A(_2473_),
    .B(\dmmu0.page_table[14][11] ),
    .C(_2463_),
    .X(_2477_));
 sky130_fd_sc_hd__a21o_1 _5299_ (.A1(_2251_),
    .A2(_2461_),
    .B1(_2477_),
    .X(_0075_));
 sky130_fd_sc_hd__and3_1 _5300_ (.A(_2473_),
    .B(\dmmu0.page_table[14][12] ),
    .C(_2463_),
    .X(_2478_));
 sky130_fd_sc_hd__a21o_1 _5301_ (.A1(_2253_),
    .A2(_2461_),
    .B1(_2478_),
    .X(_0076_));
 sky130_fd_sc_hd__or2_1 _5302_ (.A(_1922_),
    .B(_2367_),
    .X(_2479_));
 sky130_fd_sc_hd__clkbuf_4 _5303_ (.A(_2479_),
    .X(_2480_));
 sky130_fd_sc_hd__nor2_1 _5304_ (.A(_1926_),
    .B(_2479_),
    .Y(_2481_));
 sky130_fd_sc_hd__a31o_1 _5305_ (.A1(_2363_),
    .A2(\immu_0.page_table[10][0] ),
    .A3(_2480_),
    .B1(_2481_),
    .X(_0077_));
 sky130_fd_sc_hd__nor2_4 _5306_ (.A(_1930_),
    .B(_2367_),
    .Y(_2482_));
 sky130_fd_sc_hd__and2_1 _5307_ (.A(_1928_),
    .B(_2482_),
    .X(_2483_));
 sky130_fd_sc_hd__a31o_1 _5308_ (.A1(_2363_),
    .A2(\immu_0.page_table[10][1] ),
    .A3(_2480_),
    .B1(_2483_),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _5309_ (.A(_1933_),
    .B(_2482_),
    .X(_2484_));
 sky130_fd_sc_hd__a31o_1 _5310_ (.A1(_2363_),
    .A2(\immu_0.page_table[10][2] ),
    .A3(_2480_),
    .B1(_2484_),
    .X(_0079_));
 sky130_fd_sc_hd__and2_1 _5311_ (.A(_1935_),
    .B(_2482_),
    .X(_2485_));
 sky130_fd_sc_hd__a31o_1 _5312_ (.A1(_2363_),
    .A2(\immu_0.page_table[10][3] ),
    .A3(_2480_),
    .B1(_2485_),
    .X(_0080_));
 sky130_fd_sc_hd__and2_1 _5313_ (.A(_1937_),
    .B(_2482_),
    .X(_2486_));
 sky130_fd_sc_hd__a31o_1 _5314_ (.A1(_2363_),
    .A2(\immu_0.page_table[10][4] ),
    .A3(_2480_),
    .B1(_2486_),
    .X(_0081_));
 sky130_fd_sc_hd__and2_1 _5315_ (.A(_1940_),
    .B(_2482_),
    .X(_2487_));
 sky130_fd_sc_hd__a31o_1 _5316_ (.A1(_2363_),
    .A2(\immu_0.page_table[10][5] ),
    .A3(_2480_),
    .B1(_2487_),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _5317_ (.A(_1942_),
    .B(_2482_),
    .X(_2488_));
 sky130_fd_sc_hd__a31o_1 _5318_ (.A1(_2363_),
    .A2(\immu_0.page_table[10][6] ),
    .A3(_2480_),
    .B1(_2488_),
    .X(_0083_));
 sky130_fd_sc_hd__buf_4 _5319_ (.A(_2300_),
    .X(_2489_));
 sky130_fd_sc_hd__and2_1 _5320_ (.A(_1944_),
    .B(_2482_),
    .X(_2490_));
 sky130_fd_sc_hd__a31o_1 _5321_ (.A1(_2489_),
    .A2(\immu_0.page_table[10][7] ),
    .A3(_2480_),
    .B1(_2490_),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _5322_ (.A(_2310_),
    .B(_2482_),
    .X(_2491_));
 sky130_fd_sc_hd__a31o_1 _5323_ (.A1(_2489_),
    .A2(\immu_0.page_table[10][8] ),
    .A3(_2480_),
    .B1(_2491_),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _5324_ (.A(_2312_),
    .B(_2482_),
    .X(_2492_));
 sky130_fd_sc_hd__a31o_1 _5325_ (.A1(_2489_),
    .A2(\immu_0.page_table[10][9] ),
    .A3(_2480_),
    .B1(_2492_),
    .X(_0086_));
 sky130_fd_sc_hd__and2_1 _5326_ (.A(_2314_),
    .B(_2482_),
    .X(_2493_));
 sky130_fd_sc_hd__a31o_1 _5327_ (.A1(_2489_),
    .A2(\immu_0.page_table[10][10] ),
    .A3(_2479_),
    .B1(_2493_),
    .X(_0087_));
 sky130_fd_sc_hd__or2_1 _5328_ (.A(_1929_),
    .B(_2388_),
    .X(_2494_));
 sky130_fd_sc_hd__clkbuf_4 _5329_ (.A(_2494_),
    .X(_2495_));
 sky130_fd_sc_hd__nor2_1 _5330_ (.A(_1926_),
    .B(_2494_),
    .Y(_2496_));
 sky130_fd_sc_hd__a31o_1 _5331_ (.A1(_2489_),
    .A2(\immu_0.page_table[9][0] ),
    .A3(_2495_),
    .B1(_2496_),
    .X(_0088_));
 sky130_fd_sc_hd__nor2_4 _5332_ (.A(_1930_),
    .B(_2388_),
    .Y(_2497_));
 sky130_fd_sc_hd__and2_1 _5333_ (.A(_1928_),
    .B(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__a31o_1 _5334_ (.A1(_2489_),
    .A2(\immu_0.page_table[9][1] ),
    .A3(_2495_),
    .B1(_2498_),
    .X(_0089_));
 sky130_fd_sc_hd__and2_1 _5335_ (.A(_1933_),
    .B(_2497_),
    .X(_2499_));
 sky130_fd_sc_hd__a31o_1 _5336_ (.A1(_2489_),
    .A2(\immu_0.page_table[9][2] ),
    .A3(_2495_),
    .B1(_2499_),
    .X(_0090_));
 sky130_fd_sc_hd__and2_1 _5337_ (.A(_1935_),
    .B(_2497_),
    .X(_2500_));
 sky130_fd_sc_hd__a31o_1 _5338_ (.A1(_2489_),
    .A2(\immu_0.page_table[9][3] ),
    .A3(_2495_),
    .B1(_2500_),
    .X(_0091_));
 sky130_fd_sc_hd__and2_1 _5339_ (.A(_1937_),
    .B(_2497_),
    .X(_2501_));
 sky130_fd_sc_hd__a31o_1 _5340_ (.A1(_2489_),
    .A2(\immu_0.page_table[9][4] ),
    .A3(_2495_),
    .B1(_2501_),
    .X(_0092_));
 sky130_fd_sc_hd__and2_1 _5341_ (.A(_1940_),
    .B(_2497_),
    .X(_2502_));
 sky130_fd_sc_hd__a31o_1 _5342_ (.A1(_2489_),
    .A2(\immu_0.page_table[9][5] ),
    .A3(_2495_),
    .B1(_2502_),
    .X(_0093_));
 sky130_fd_sc_hd__clkbuf_4 _5343_ (.A(_2300_),
    .X(_2503_));
 sky130_fd_sc_hd__and2_1 _5344_ (.A(_1942_),
    .B(_2497_),
    .X(_2504_));
 sky130_fd_sc_hd__a31o_1 _5345_ (.A1(_2503_),
    .A2(\immu_0.page_table[9][6] ),
    .A3(_2495_),
    .B1(_2504_),
    .X(_0094_));
 sky130_fd_sc_hd__and2_1 _5346_ (.A(_1944_),
    .B(_2497_),
    .X(_2505_));
 sky130_fd_sc_hd__a31o_1 _5347_ (.A1(_2503_),
    .A2(\immu_0.page_table[9][7] ),
    .A3(_2495_),
    .B1(_2505_),
    .X(_0095_));
 sky130_fd_sc_hd__and2_1 _5348_ (.A(_2310_),
    .B(_2497_),
    .X(_2506_));
 sky130_fd_sc_hd__a31o_1 _5349_ (.A1(_2503_),
    .A2(\immu_0.page_table[9][8] ),
    .A3(_2495_),
    .B1(_2506_),
    .X(_0096_));
 sky130_fd_sc_hd__and2_1 _5350_ (.A(_2312_),
    .B(_2497_),
    .X(_2507_));
 sky130_fd_sc_hd__a31o_1 _5351_ (.A1(_2503_),
    .A2(\immu_0.page_table[9][9] ),
    .A3(_2495_),
    .B1(_2507_),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _5352_ (.A(_2314_),
    .B(_2497_),
    .X(_2508_));
 sky130_fd_sc_hd__a31o_1 _5353_ (.A1(_2503_),
    .A2(\immu_0.page_table[9][10] ),
    .A3(_2494_),
    .B1(_2508_),
    .X(_0098_));
 sky130_fd_sc_hd__or2_1 _5354_ (.A(_1929_),
    .B(_2407_),
    .X(_2509_));
 sky130_fd_sc_hd__clkbuf_4 _5355_ (.A(_2509_),
    .X(_2510_));
 sky130_fd_sc_hd__nor2_1 _5356_ (.A(_1926_),
    .B(_2509_),
    .Y(_2511_));
 sky130_fd_sc_hd__a31o_1 _5357_ (.A1(_2503_),
    .A2(\immu_0.page_table[8][0] ),
    .A3(_2510_),
    .B1(_2511_),
    .X(_0099_));
 sky130_fd_sc_hd__nor2_4 _5358_ (.A(_1930_),
    .B(_2407_),
    .Y(_2512_));
 sky130_fd_sc_hd__and2_1 _5359_ (.A(_1928_),
    .B(_2512_),
    .X(_2513_));
 sky130_fd_sc_hd__a31o_1 _5360_ (.A1(_2503_),
    .A2(\immu_0.page_table[8][1] ),
    .A3(_2510_),
    .B1(_2513_),
    .X(_0100_));
 sky130_fd_sc_hd__and2_1 _5361_ (.A(_1933_),
    .B(_2512_),
    .X(_2514_));
 sky130_fd_sc_hd__a31o_1 _5362_ (.A1(_2503_),
    .A2(\immu_0.page_table[8][2] ),
    .A3(_2510_),
    .B1(_2514_),
    .X(_0101_));
 sky130_fd_sc_hd__and2_1 _5363_ (.A(_1935_),
    .B(_2512_),
    .X(_2515_));
 sky130_fd_sc_hd__a31o_1 _5364_ (.A1(_2503_),
    .A2(\immu_0.page_table[8][3] ),
    .A3(_2510_),
    .B1(_2515_),
    .X(_0102_));
 sky130_fd_sc_hd__and2_1 _5365_ (.A(_1937_),
    .B(_2512_),
    .X(_2516_));
 sky130_fd_sc_hd__a31o_1 _5366_ (.A1(_2503_),
    .A2(\immu_0.page_table[8][4] ),
    .A3(_2510_),
    .B1(_2516_),
    .X(_0103_));
 sky130_fd_sc_hd__clkbuf_4 _5367_ (.A(_2300_),
    .X(_2517_));
 sky130_fd_sc_hd__and2_1 _5368_ (.A(_1940_),
    .B(_2512_),
    .X(_2518_));
 sky130_fd_sc_hd__a31o_1 _5369_ (.A1(_2517_),
    .A2(\immu_0.page_table[8][5] ),
    .A3(_2510_),
    .B1(_2518_),
    .X(_0104_));
 sky130_fd_sc_hd__and2_1 _5370_ (.A(_1942_),
    .B(_2512_),
    .X(_2519_));
 sky130_fd_sc_hd__a31o_1 _5371_ (.A1(_2517_),
    .A2(\immu_0.page_table[8][6] ),
    .A3(_2510_),
    .B1(_2519_),
    .X(_0105_));
 sky130_fd_sc_hd__and2_1 _5372_ (.A(_1944_),
    .B(_2512_),
    .X(_2520_));
 sky130_fd_sc_hd__a31o_1 _5373_ (.A1(_2517_),
    .A2(\immu_0.page_table[8][7] ),
    .A3(_2510_),
    .B1(_2520_),
    .X(_0106_));
 sky130_fd_sc_hd__and2_1 _5374_ (.A(_2310_),
    .B(_2512_),
    .X(_2521_));
 sky130_fd_sc_hd__a31o_1 _5375_ (.A1(_2517_),
    .A2(\immu_0.page_table[8][8] ),
    .A3(_2510_),
    .B1(_2521_),
    .X(_0107_));
 sky130_fd_sc_hd__and2_1 _5376_ (.A(_2312_),
    .B(_2512_),
    .X(_2522_));
 sky130_fd_sc_hd__a31o_1 _5377_ (.A1(_2517_),
    .A2(\immu_0.page_table[8][9] ),
    .A3(_2510_),
    .B1(_2522_),
    .X(_0108_));
 sky130_fd_sc_hd__and2_1 _5378_ (.A(_2314_),
    .B(_2512_),
    .X(_2523_));
 sky130_fd_sc_hd__a31o_1 _5379_ (.A1(_2517_),
    .A2(\immu_0.page_table[8][10] ),
    .A3(_2509_),
    .B1(_2523_),
    .X(_0109_));
 sky130_fd_sc_hd__or2_1 _5380_ (.A(_1929_),
    .B(_2440_),
    .X(_2524_));
 sky130_fd_sc_hd__clkbuf_4 _5381_ (.A(_2524_),
    .X(_2525_));
 sky130_fd_sc_hd__nor2_1 _5382_ (.A(_1926_),
    .B(_2524_),
    .Y(_2526_));
 sky130_fd_sc_hd__a31o_1 _5383_ (.A1(_2517_),
    .A2(\immu_0.page_table[7][0] ),
    .A3(_2525_),
    .B1(_2526_),
    .X(_0110_));
 sky130_fd_sc_hd__nor2_4 _5384_ (.A(_1930_),
    .B(_2440_),
    .Y(_2527_));
 sky130_fd_sc_hd__and2_1 _5385_ (.A(net96),
    .B(_2527_),
    .X(_2528_));
 sky130_fd_sc_hd__a31o_1 _5386_ (.A1(_2517_),
    .A2(\immu_0.page_table[7][1] ),
    .A3(_2525_),
    .B1(_2528_),
    .X(_0111_));
 sky130_fd_sc_hd__and2_1 _5387_ (.A(_1933_),
    .B(_2527_),
    .X(_2529_));
 sky130_fd_sc_hd__a31o_1 _5388_ (.A1(_2517_),
    .A2(\immu_0.page_table[7][2] ),
    .A3(_2525_),
    .B1(_2529_),
    .X(_0112_));
 sky130_fd_sc_hd__and2_1 _5389_ (.A(_1935_),
    .B(_2527_),
    .X(_2530_));
 sky130_fd_sc_hd__a31o_1 _5390_ (.A1(_2517_),
    .A2(\immu_0.page_table[7][3] ),
    .A3(_2525_),
    .B1(_2530_),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_4 _5391_ (.A(_2300_),
    .X(_2531_));
 sky130_fd_sc_hd__and2_1 _5392_ (.A(_1937_),
    .B(_2527_),
    .X(_2532_));
 sky130_fd_sc_hd__a31o_1 _5393_ (.A1(_2531_),
    .A2(\immu_0.page_table[7][4] ),
    .A3(_2525_),
    .B1(_2532_),
    .X(_0114_));
 sky130_fd_sc_hd__and2_1 _5394_ (.A(_1940_),
    .B(_2527_),
    .X(_2533_));
 sky130_fd_sc_hd__a31o_1 _5395_ (.A1(_2531_),
    .A2(\immu_0.page_table[7][5] ),
    .A3(_2525_),
    .B1(_2533_),
    .X(_0115_));
 sky130_fd_sc_hd__and2_1 _5396_ (.A(_1942_),
    .B(_2527_),
    .X(_2534_));
 sky130_fd_sc_hd__a31o_1 _5397_ (.A1(_2531_),
    .A2(\immu_0.page_table[7][6] ),
    .A3(_2525_),
    .B1(_2534_),
    .X(_0116_));
 sky130_fd_sc_hd__and2_1 _5398_ (.A(_1944_),
    .B(_2527_),
    .X(_2535_));
 sky130_fd_sc_hd__a31o_1 _5399_ (.A1(_2531_),
    .A2(\immu_0.page_table[7][7] ),
    .A3(_2525_),
    .B1(_2535_),
    .X(_0117_));
 sky130_fd_sc_hd__and2_1 _5400_ (.A(_2310_),
    .B(_2527_),
    .X(_2536_));
 sky130_fd_sc_hd__a31o_1 _5401_ (.A1(_2531_),
    .A2(\immu_0.page_table[7][8] ),
    .A3(_2525_),
    .B1(_2536_),
    .X(_0118_));
 sky130_fd_sc_hd__and2_1 _5402_ (.A(_2312_),
    .B(_2527_),
    .X(_2537_));
 sky130_fd_sc_hd__a31o_1 _5403_ (.A1(_2531_),
    .A2(\immu_0.page_table[7][9] ),
    .A3(_2525_),
    .B1(_2537_),
    .X(_0119_));
 sky130_fd_sc_hd__and2_1 _5404_ (.A(_2314_),
    .B(_2527_),
    .X(_2538_));
 sky130_fd_sc_hd__a31o_1 _5405_ (.A1(_2531_),
    .A2(\immu_0.page_table[7][10] ),
    .A3(_2524_),
    .B1(_2538_),
    .X(_0120_));
 sky130_fd_sc_hd__or2_4 _5406_ (.A(_2317_),
    .B(_2439_),
    .X(_2539_));
 sky130_fd_sc_hd__or2_1 _5407_ (.A(_1929_),
    .B(_2539_),
    .X(_2540_));
 sky130_fd_sc_hd__clkbuf_4 _5408_ (.A(_2540_),
    .X(_2541_));
 sky130_fd_sc_hd__nor2_1 _5409_ (.A(_1925_),
    .B(_2540_),
    .Y(_2542_));
 sky130_fd_sc_hd__a31o_1 _5410_ (.A1(_2531_),
    .A2(\immu_0.page_table[6][0] ),
    .A3(_2541_),
    .B1(_2542_),
    .X(_0121_));
 sky130_fd_sc_hd__nor2_4 _5411_ (.A(_1930_),
    .B(_2539_),
    .Y(_2543_));
 sky130_fd_sc_hd__and2_1 _5412_ (.A(net96),
    .B(_2543_),
    .X(_2544_));
 sky130_fd_sc_hd__a31o_1 _5413_ (.A1(_2531_),
    .A2(\immu_0.page_table[6][1] ),
    .A3(_2541_),
    .B1(_2544_),
    .X(_0122_));
 sky130_fd_sc_hd__and2_1 _5414_ (.A(net97),
    .B(_2543_),
    .X(_2545_));
 sky130_fd_sc_hd__a31o_1 _5415_ (.A1(_2531_),
    .A2(\immu_0.page_table[6][2] ),
    .A3(_2541_),
    .B1(_2545_),
    .X(_0123_));
 sky130_fd_sc_hd__clkbuf_4 _5416_ (.A(_2300_),
    .X(_2546_));
 sky130_fd_sc_hd__and2_1 _5417_ (.A(net98),
    .B(_2543_),
    .X(_2547_));
 sky130_fd_sc_hd__a31o_1 _5418_ (.A1(_2546_),
    .A2(\immu_0.page_table[6][3] ),
    .A3(_2541_),
    .B1(_2547_),
    .X(_0124_));
 sky130_fd_sc_hd__and2_1 _5419_ (.A(net99),
    .B(_2543_),
    .X(_2548_));
 sky130_fd_sc_hd__a31o_1 _5420_ (.A1(_2546_),
    .A2(\immu_0.page_table[6][4] ),
    .A3(_2541_),
    .B1(_2548_),
    .X(_0125_));
 sky130_fd_sc_hd__and2_1 _5421_ (.A(net100),
    .B(_2543_),
    .X(_2549_));
 sky130_fd_sc_hd__a31o_1 _5422_ (.A1(_2546_),
    .A2(\immu_0.page_table[6][5] ),
    .A3(_2541_),
    .B1(_2549_),
    .X(_0126_));
 sky130_fd_sc_hd__and2_1 _5423_ (.A(net101),
    .B(_2543_),
    .X(_2550_));
 sky130_fd_sc_hd__a31o_1 _5424_ (.A1(_2546_),
    .A2(\immu_0.page_table[6][6] ),
    .A3(_2541_),
    .B1(_2550_),
    .X(_0127_));
 sky130_fd_sc_hd__and2_1 _5425_ (.A(net102),
    .B(_2543_),
    .X(_2551_));
 sky130_fd_sc_hd__a31o_1 _5426_ (.A1(_2546_),
    .A2(\immu_0.page_table[6][7] ),
    .A3(_2541_),
    .B1(_2551_),
    .X(_0128_));
 sky130_fd_sc_hd__and2_1 _5427_ (.A(_2310_),
    .B(_2543_),
    .X(_2552_));
 sky130_fd_sc_hd__a31o_1 _5428_ (.A1(_2546_),
    .A2(\immu_0.page_table[6][8] ),
    .A3(_2541_),
    .B1(_2552_),
    .X(_0129_));
 sky130_fd_sc_hd__and2_1 _5429_ (.A(_2312_),
    .B(_2543_),
    .X(_2553_));
 sky130_fd_sc_hd__a31o_1 _5430_ (.A1(_2546_),
    .A2(\immu_0.page_table[6][9] ),
    .A3(_2541_),
    .B1(_2553_),
    .X(_0130_));
 sky130_fd_sc_hd__and2_1 _5431_ (.A(_2314_),
    .B(_2543_),
    .X(_2554_));
 sky130_fd_sc_hd__a31o_1 _5432_ (.A1(_2546_),
    .A2(\immu_0.page_table[6][10] ),
    .A3(_2540_),
    .B1(_2554_),
    .X(_0131_));
 sky130_fd_sc_hd__or2_4 _5433_ (.A(_2350_),
    .B(_2439_),
    .X(_2555_));
 sky130_fd_sc_hd__or2_1 _5434_ (.A(_1929_),
    .B(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__clkbuf_4 _5435_ (.A(_2556_),
    .X(_2557_));
 sky130_fd_sc_hd__nor2_1 _5436_ (.A(_1925_),
    .B(_2556_),
    .Y(_2558_));
 sky130_fd_sc_hd__a31o_1 _5437_ (.A1(_2546_),
    .A2(\immu_0.page_table[5][0] ),
    .A3(_2557_),
    .B1(_2558_),
    .X(_0132_));
 sky130_fd_sc_hd__nor2_4 _5438_ (.A(_1922_),
    .B(_2555_),
    .Y(_2559_));
 sky130_fd_sc_hd__and2_1 _5439_ (.A(net96),
    .B(_2559_),
    .X(_2560_));
 sky130_fd_sc_hd__a31o_1 _5440_ (.A1(_2546_),
    .A2(\immu_0.page_table[5][1] ),
    .A3(_2557_),
    .B1(_2560_),
    .X(_0133_));
 sky130_fd_sc_hd__buf_4 _5441_ (.A(_1897_),
    .X(_2561_));
 sky130_fd_sc_hd__clkbuf_4 _5442_ (.A(_2561_),
    .X(_2562_));
 sky130_fd_sc_hd__and2_1 _5443_ (.A(net97),
    .B(_2559_),
    .X(_2563_));
 sky130_fd_sc_hd__a31o_1 _5444_ (.A1(_2562_),
    .A2(\immu_0.page_table[5][2] ),
    .A3(_2557_),
    .B1(_2563_),
    .X(_0134_));
 sky130_fd_sc_hd__and2_1 _5445_ (.A(net98),
    .B(_2559_),
    .X(_2564_));
 sky130_fd_sc_hd__a31o_1 _5446_ (.A1(_2562_),
    .A2(\immu_0.page_table[5][3] ),
    .A3(_2557_),
    .B1(_2564_),
    .X(_0135_));
 sky130_fd_sc_hd__and2_1 _5447_ (.A(net99),
    .B(_2559_),
    .X(_2565_));
 sky130_fd_sc_hd__a31o_1 _5448_ (.A1(_2562_),
    .A2(\immu_0.page_table[5][4] ),
    .A3(_2557_),
    .B1(_2565_),
    .X(_0136_));
 sky130_fd_sc_hd__and2_1 _5449_ (.A(net100),
    .B(_2559_),
    .X(_2566_));
 sky130_fd_sc_hd__a31o_1 _5450_ (.A1(_2562_),
    .A2(\immu_0.page_table[5][5] ),
    .A3(_2557_),
    .B1(_2566_),
    .X(_0137_));
 sky130_fd_sc_hd__and2_1 _5451_ (.A(net101),
    .B(_2559_),
    .X(_2567_));
 sky130_fd_sc_hd__a31o_1 _5452_ (.A1(_2562_),
    .A2(\immu_0.page_table[5][6] ),
    .A3(_2557_),
    .B1(_2567_),
    .X(_0138_));
 sky130_fd_sc_hd__and2_1 _5453_ (.A(net102),
    .B(_2559_),
    .X(_2568_));
 sky130_fd_sc_hd__a31o_1 _5454_ (.A1(_2562_),
    .A2(\immu_0.page_table[5][7] ),
    .A3(_2557_),
    .B1(_2568_),
    .X(_0139_));
 sky130_fd_sc_hd__and2_1 _5455_ (.A(_2310_),
    .B(_2559_),
    .X(_2569_));
 sky130_fd_sc_hd__a31o_1 _5456_ (.A1(_2562_),
    .A2(\immu_0.page_table[5][8] ),
    .A3(_2557_),
    .B1(_2569_),
    .X(_0140_));
 sky130_fd_sc_hd__and2_1 _5457_ (.A(_2312_),
    .B(_2559_),
    .X(_2570_));
 sky130_fd_sc_hd__a31o_1 _5458_ (.A1(_2562_),
    .A2(\immu_0.page_table[5][9] ),
    .A3(_2557_),
    .B1(_2570_),
    .X(_0141_));
 sky130_fd_sc_hd__and2_1 _5459_ (.A(_2314_),
    .B(_2559_),
    .X(_2571_));
 sky130_fd_sc_hd__a31o_1 _5460_ (.A1(_2562_),
    .A2(\immu_0.page_table[5][10] ),
    .A3(_2556_),
    .B1(_2571_),
    .X(_0142_));
 sky130_fd_sc_hd__or3_4 _5461_ (.A(net83),
    .B(net76),
    .C(_2439_),
    .X(_2572_));
 sky130_fd_sc_hd__or2_1 _5462_ (.A(_1929_),
    .B(_2572_),
    .X(_2573_));
 sky130_fd_sc_hd__clkbuf_4 _5463_ (.A(_2573_),
    .X(_2574_));
 sky130_fd_sc_hd__nor2_1 _5464_ (.A(_1925_),
    .B(_2573_),
    .Y(_2575_));
 sky130_fd_sc_hd__a31o_1 _5465_ (.A1(_2562_),
    .A2(\immu_0.page_table[4][0] ),
    .A3(_2574_),
    .B1(_2575_),
    .X(_0143_));
 sky130_fd_sc_hd__clkbuf_4 _5466_ (.A(_2561_),
    .X(_2576_));
 sky130_fd_sc_hd__nor2_4 _5467_ (.A(_1922_),
    .B(_2572_),
    .Y(_2577_));
 sky130_fd_sc_hd__and2_1 _5468_ (.A(net96),
    .B(_2577_),
    .X(_2578_));
 sky130_fd_sc_hd__a31o_1 _5469_ (.A1(_2576_),
    .A2(\immu_0.page_table[4][1] ),
    .A3(_2574_),
    .B1(_2578_),
    .X(_0144_));
 sky130_fd_sc_hd__and2_1 _5470_ (.A(net97),
    .B(_2577_),
    .X(_2579_));
 sky130_fd_sc_hd__a31o_1 _5471_ (.A1(_2576_),
    .A2(\immu_0.page_table[4][2] ),
    .A3(_2574_),
    .B1(_2579_),
    .X(_0145_));
 sky130_fd_sc_hd__and2_1 _5472_ (.A(net98),
    .B(_2577_),
    .X(_2580_));
 sky130_fd_sc_hd__a31o_1 _5473_ (.A1(_2576_),
    .A2(\immu_0.page_table[4][3] ),
    .A3(_2574_),
    .B1(_2580_),
    .X(_0146_));
 sky130_fd_sc_hd__and2_1 _5474_ (.A(net99),
    .B(_2577_),
    .X(_2581_));
 sky130_fd_sc_hd__a31o_1 _5475_ (.A1(_2576_),
    .A2(\immu_0.page_table[4][4] ),
    .A3(_2574_),
    .B1(_2581_),
    .X(_0147_));
 sky130_fd_sc_hd__and2_1 _5476_ (.A(net100),
    .B(_2577_),
    .X(_2582_));
 sky130_fd_sc_hd__a31o_1 _5477_ (.A1(_2576_),
    .A2(\immu_0.page_table[4][5] ),
    .A3(_2574_),
    .B1(_2582_),
    .X(_0148_));
 sky130_fd_sc_hd__and2_1 _5478_ (.A(net101),
    .B(_2577_),
    .X(_2583_));
 sky130_fd_sc_hd__a31o_1 _5479_ (.A1(_2576_),
    .A2(\immu_0.page_table[4][6] ),
    .A3(_2574_),
    .B1(_2583_),
    .X(_0149_));
 sky130_fd_sc_hd__and2_1 _5480_ (.A(net102),
    .B(_2577_),
    .X(_2584_));
 sky130_fd_sc_hd__a31o_1 _5481_ (.A1(_2576_),
    .A2(\immu_0.page_table[4][7] ),
    .A3(_2574_),
    .B1(_2584_),
    .X(_0150_));
 sky130_fd_sc_hd__and2_1 _5482_ (.A(net103),
    .B(_2577_),
    .X(_2585_));
 sky130_fd_sc_hd__a31o_1 _5483_ (.A1(_2576_),
    .A2(\immu_0.page_table[4][8] ),
    .A3(_2574_),
    .B1(_2585_),
    .X(_0151_));
 sky130_fd_sc_hd__and2_1 _5484_ (.A(net104),
    .B(_2577_),
    .X(_2586_));
 sky130_fd_sc_hd__a31o_1 _5485_ (.A1(_2576_),
    .A2(\immu_0.page_table[4][9] ),
    .A3(_2574_),
    .B1(_2586_),
    .X(_0152_));
 sky130_fd_sc_hd__and2_1 _5486_ (.A(net93),
    .B(_2577_),
    .X(_2587_));
 sky130_fd_sc_hd__a31o_1 _5487_ (.A1(_2576_),
    .A2(\immu_0.page_table[4][10] ),
    .A3(_2573_),
    .B1(_2587_),
    .X(_0153_));
 sky130_fd_sc_hd__clkbuf_4 _5488_ (.A(_2561_),
    .X(_2588_));
 sky130_fd_sc_hd__or3_4 _5489_ (.A(net85),
    .B(net84),
    .C(_1912_),
    .X(_2589_));
 sky130_fd_sc_hd__or2_1 _5490_ (.A(_1929_),
    .B(_2589_),
    .X(_2590_));
 sky130_fd_sc_hd__clkbuf_4 _5491_ (.A(_2590_),
    .X(_2591_));
 sky130_fd_sc_hd__nor2_1 _5492_ (.A(_1925_),
    .B(_2590_),
    .Y(_2592_));
 sky130_fd_sc_hd__a31o_1 _5493_ (.A1(_2588_),
    .A2(\immu_0.page_table[3][0] ),
    .A3(_2591_),
    .B1(_2592_),
    .X(_0154_));
 sky130_fd_sc_hd__nor2_4 _5494_ (.A(_1922_),
    .B(_2589_),
    .Y(_2593_));
 sky130_fd_sc_hd__and2_1 _5495_ (.A(net96),
    .B(_2593_),
    .X(_2594_));
 sky130_fd_sc_hd__a31o_1 _5496_ (.A1(_2588_),
    .A2(\immu_0.page_table[3][1] ),
    .A3(_2591_),
    .B1(_2594_),
    .X(_0155_));
 sky130_fd_sc_hd__and2_1 _5497_ (.A(net97),
    .B(_2593_),
    .X(_2595_));
 sky130_fd_sc_hd__a31o_1 _5498_ (.A1(_2588_),
    .A2(\immu_0.page_table[3][2] ),
    .A3(_2591_),
    .B1(_2595_),
    .X(_0156_));
 sky130_fd_sc_hd__and2_1 _5499_ (.A(net98),
    .B(_2593_),
    .X(_2596_));
 sky130_fd_sc_hd__a31o_1 _5500_ (.A1(_2588_),
    .A2(\immu_0.page_table[3][3] ),
    .A3(_2591_),
    .B1(_2596_),
    .X(_0157_));
 sky130_fd_sc_hd__and2_1 _5501_ (.A(net99),
    .B(_2593_),
    .X(_2597_));
 sky130_fd_sc_hd__a31o_1 _5502_ (.A1(_2588_),
    .A2(\immu_0.page_table[3][4] ),
    .A3(_2591_),
    .B1(_2597_),
    .X(_0158_));
 sky130_fd_sc_hd__and2_1 _5503_ (.A(net100),
    .B(_2593_),
    .X(_2598_));
 sky130_fd_sc_hd__a31o_1 _5504_ (.A1(_2588_),
    .A2(\immu_0.page_table[3][5] ),
    .A3(_2591_),
    .B1(_2598_),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _5505_ (.A(net101),
    .B(_2593_),
    .X(_2599_));
 sky130_fd_sc_hd__a31o_1 _5506_ (.A1(_2588_),
    .A2(\immu_0.page_table[3][6] ),
    .A3(_2591_),
    .B1(_2599_),
    .X(_0160_));
 sky130_fd_sc_hd__and2_1 _5507_ (.A(net102),
    .B(_2593_),
    .X(_2600_));
 sky130_fd_sc_hd__a31o_1 _5508_ (.A1(_2588_),
    .A2(\immu_0.page_table[3][7] ),
    .A3(_2591_),
    .B1(_2600_),
    .X(_0161_));
 sky130_fd_sc_hd__and2_1 _5509_ (.A(net103),
    .B(_2593_),
    .X(_2601_));
 sky130_fd_sc_hd__a31o_1 _5510_ (.A1(_2588_),
    .A2(\immu_0.page_table[3][8] ),
    .A3(_2591_),
    .B1(_2601_),
    .X(_0162_));
 sky130_fd_sc_hd__and2_1 _5511_ (.A(net104),
    .B(_2593_),
    .X(_2602_));
 sky130_fd_sc_hd__a31o_1 _5512_ (.A1(_2588_),
    .A2(\immu_0.page_table[3][9] ),
    .A3(_2591_),
    .B1(_2602_),
    .X(_0163_));
 sky130_fd_sc_hd__clkbuf_4 _5513_ (.A(_2561_),
    .X(_2603_));
 sky130_fd_sc_hd__and2_1 _5514_ (.A(net93),
    .B(_2593_),
    .X(_2604_));
 sky130_fd_sc_hd__a31o_1 _5515_ (.A1(_2603_),
    .A2(\immu_0.page_table[3][10] ),
    .A3(_2590_),
    .B1(_2604_),
    .X(_0164_));
 sky130_fd_sc_hd__or3_4 _5516_ (.A(net85),
    .B(net84),
    .C(_2317_),
    .X(_2605_));
 sky130_fd_sc_hd__or2_1 _5517_ (.A(_1929_),
    .B(_2605_),
    .X(_2606_));
 sky130_fd_sc_hd__clkbuf_4 _5518_ (.A(_2606_),
    .X(_2607_));
 sky130_fd_sc_hd__nor2_1 _5519_ (.A(_1925_),
    .B(_2606_),
    .Y(_2608_));
 sky130_fd_sc_hd__a31o_1 _5520_ (.A1(_2603_),
    .A2(\immu_0.page_table[2][0] ),
    .A3(_2607_),
    .B1(_2608_),
    .X(_0165_));
 sky130_fd_sc_hd__nor2_4 _5521_ (.A(_1922_),
    .B(_2605_),
    .Y(_2609_));
 sky130_fd_sc_hd__and2_1 _5522_ (.A(net96),
    .B(_2609_),
    .X(_2610_));
 sky130_fd_sc_hd__a31o_1 _5523_ (.A1(_2603_),
    .A2(\immu_0.page_table[2][1] ),
    .A3(_2607_),
    .B1(_2610_),
    .X(_0166_));
 sky130_fd_sc_hd__and2_1 _5524_ (.A(net97),
    .B(_2609_),
    .X(_2611_));
 sky130_fd_sc_hd__a31o_1 _5525_ (.A1(_2603_),
    .A2(\immu_0.page_table[2][2] ),
    .A3(_2607_),
    .B1(_2611_),
    .X(_0167_));
 sky130_fd_sc_hd__and2_1 _5526_ (.A(net98),
    .B(_2609_),
    .X(_2612_));
 sky130_fd_sc_hd__a31o_1 _5527_ (.A1(_2603_),
    .A2(\immu_0.page_table[2][3] ),
    .A3(_2607_),
    .B1(_2612_),
    .X(_0168_));
 sky130_fd_sc_hd__and2_1 _5528_ (.A(net99),
    .B(_2609_),
    .X(_2613_));
 sky130_fd_sc_hd__a31o_1 _5529_ (.A1(_2603_),
    .A2(\immu_0.page_table[2][4] ),
    .A3(_2607_),
    .B1(_2613_),
    .X(_0169_));
 sky130_fd_sc_hd__and2_1 _5530_ (.A(net100),
    .B(_2609_),
    .X(_2614_));
 sky130_fd_sc_hd__a31o_1 _5531_ (.A1(_2603_),
    .A2(\immu_0.page_table[2][5] ),
    .A3(_2607_),
    .B1(_2614_),
    .X(_0170_));
 sky130_fd_sc_hd__and2_1 _5532_ (.A(net101),
    .B(_2609_),
    .X(_2615_));
 sky130_fd_sc_hd__a31o_1 _5533_ (.A1(_2603_),
    .A2(\immu_0.page_table[2][6] ),
    .A3(_2607_),
    .B1(_2615_),
    .X(_0171_));
 sky130_fd_sc_hd__and2_1 _5534_ (.A(net102),
    .B(_2609_),
    .X(_2616_));
 sky130_fd_sc_hd__a31o_1 _5535_ (.A1(_2603_),
    .A2(\immu_0.page_table[2][7] ),
    .A3(_2607_),
    .B1(_2616_),
    .X(_0172_));
 sky130_fd_sc_hd__and2_1 _5536_ (.A(net103),
    .B(_2609_),
    .X(_2617_));
 sky130_fd_sc_hd__a31o_1 _5537_ (.A1(_2603_),
    .A2(\immu_0.page_table[2][8] ),
    .A3(_2607_),
    .B1(_2617_),
    .X(_0173_));
 sky130_fd_sc_hd__buf_4 _5538_ (.A(_2561_),
    .X(_2618_));
 sky130_fd_sc_hd__and2_1 _5539_ (.A(net104),
    .B(_2609_),
    .X(_2619_));
 sky130_fd_sc_hd__a31o_1 _5540_ (.A1(_2618_),
    .A2(\immu_0.page_table[2][9] ),
    .A3(_2607_),
    .B1(_2619_),
    .X(_0174_));
 sky130_fd_sc_hd__and2_1 _5541_ (.A(net93),
    .B(_2609_),
    .X(_2620_));
 sky130_fd_sc_hd__a31o_1 _5542_ (.A1(_2618_),
    .A2(\immu_0.page_table[2][10] ),
    .A3(_2606_),
    .B1(_2620_),
    .X(_0175_));
 sky130_fd_sc_hd__or3_4 _5543_ (.A(net85),
    .B(net84),
    .C(_2350_),
    .X(_2621_));
 sky130_fd_sc_hd__or2_1 _5544_ (.A(_1921_),
    .B(_2621_),
    .X(_2622_));
 sky130_fd_sc_hd__clkbuf_4 _5545_ (.A(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__nand2_1 _5546_ (.A(_2190_),
    .B(_2622_),
    .Y(_2624_));
 sky130_fd_sc_hd__clkbuf_4 _5547_ (.A(_2624_),
    .X(_2625_));
 sky130_fd_sc_hd__o22a_1 _5548_ (.A1(_2210_),
    .A2(_2623_),
    .B1(_2625_),
    .B2(\immu_0.page_table[1][0] ),
    .X(_0176_));
 sky130_fd_sc_hd__o22a_1 _5549_ (.A1(_2223_),
    .A2(_2623_),
    .B1(_2625_),
    .B2(\immu_0.page_table[1][1] ),
    .X(_0177_));
 sky130_fd_sc_hd__o22a_1 _5550_ (.A1(_2226_),
    .A2(_2623_),
    .B1(_2625_),
    .B2(\immu_0.page_table[1][2] ),
    .X(_0178_));
 sky130_fd_sc_hd__o22a_1 _5551_ (.A1(_2229_),
    .A2(_2623_),
    .B1(_2625_),
    .B2(\immu_0.page_table[1][3] ),
    .X(_0179_));
 sky130_fd_sc_hd__o22a_1 _5552_ (.A1(_2232_),
    .A2(_2623_),
    .B1(_2625_),
    .B2(\immu_0.page_table[1][4] ),
    .X(_0180_));
 sky130_fd_sc_hd__o22a_1 _5553_ (.A1(_2235_),
    .A2(_2623_),
    .B1(_2625_),
    .B2(\immu_0.page_table[1][5] ),
    .X(_0181_));
 sky130_fd_sc_hd__o22a_1 _5554_ (.A1(_2239_),
    .A2(_2623_),
    .B1(_2625_),
    .B2(\immu_0.page_table[1][6] ),
    .X(_0182_));
 sky130_fd_sc_hd__o22a_1 _5555_ (.A1(_2242_),
    .A2(_2623_),
    .B1(_2625_),
    .B2(\immu_0.page_table[1][7] ),
    .X(_0183_));
 sky130_fd_sc_hd__o22a_1 _5556_ (.A1(_1946_),
    .A2(_2623_),
    .B1(_2625_),
    .B2(\immu_0.page_table[1][8] ),
    .X(_0184_));
 sky130_fd_sc_hd__o22a_1 _5557_ (.A1(_1948_),
    .A2(_2623_),
    .B1(_2625_),
    .B2(\immu_0.page_table[1][9] ),
    .X(_0185_));
 sky130_fd_sc_hd__o22a_1 _5558_ (.A1(_1950_),
    .A2(_2622_),
    .B1(_2624_),
    .B2(\immu_0.page_table[1][10] ),
    .X(_0186_));
 sky130_fd_sc_hd__or2_1 _5559_ (.A(_1929_),
    .B(_2212_),
    .X(_2626_));
 sky130_fd_sc_hd__clkbuf_4 _5560_ (.A(_2626_),
    .X(_2627_));
 sky130_fd_sc_hd__nand2_1 _5561_ (.A(_2190_),
    .B(_2626_),
    .Y(_2628_));
 sky130_fd_sc_hd__inv_2 _5562_ (.A(_2628_),
    .Y(_2629_));
 sky130_fd_sc_hd__a2bb2o_1 _5563_ (.A1_N(_1926_),
    .A2_N(_2627_),
    .B1(_2629_),
    .B2(\immu_0.page_table[0][0] ),
    .X(_0187_));
 sky130_fd_sc_hd__clkbuf_4 _5564_ (.A(_2628_),
    .X(_2630_));
 sky130_fd_sc_hd__o22a_1 _5565_ (.A1(_2223_),
    .A2(_2627_),
    .B1(_2630_),
    .B2(\immu_0.page_table[0][1] ),
    .X(_0188_));
 sky130_fd_sc_hd__o22a_1 _5566_ (.A1(_2226_),
    .A2(_2627_),
    .B1(_2630_),
    .B2(\immu_0.page_table[0][2] ),
    .X(_0189_));
 sky130_fd_sc_hd__o22a_1 _5567_ (.A1(_2229_),
    .A2(_2627_),
    .B1(_2630_),
    .B2(\immu_0.page_table[0][3] ),
    .X(_0190_));
 sky130_fd_sc_hd__o22a_1 _5568_ (.A1(_2232_),
    .A2(_2627_),
    .B1(_2630_),
    .B2(\immu_0.page_table[0][4] ),
    .X(_0191_));
 sky130_fd_sc_hd__o22a_1 _5569_ (.A1(_2235_),
    .A2(_2627_),
    .B1(_2630_),
    .B2(\immu_0.page_table[0][5] ),
    .X(_0192_));
 sky130_fd_sc_hd__o22a_1 _5570_ (.A1(_2239_),
    .A2(_2627_),
    .B1(_2630_),
    .B2(\immu_0.page_table[0][6] ),
    .X(_0193_));
 sky130_fd_sc_hd__o22a_1 _5571_ (.A1(_2242_),
    .A2(_2627_),
    .B1(_2630_),
    .B2(\immu_0.page_table[0][7] ),
    .X(_0194_));
 sky130_fd_sc_hd__o22a_1 _5572_ (.A1(_1946_),
    .A2(_2627_),
    .B1(_2630_),
    .B2(\immu_0.page_table[0][8] ),
    .X(_0195_));
 sky130_fd_sc_hd__o22a_1 _5573_ (.A1(_1948_),
    .A2(_2627_),
    .B1(_2630_),
    .B2(\immu_0.page_table[0][9] ),
    .X(_0196_));
 sky130_fd_sc_hd__o22a_1 _5574_ (.A1(_1950_),
    .A2(_2626_),
    .B1(_2630_),
    .B2(\immu_0.page_table[0][10] ),
    .X(_0197_));
 sky130_fd_sc_hd__nor2_2 _5575_ (.A(_2217_),
    .B(_2334_),
    .Y(_2631_));
 sky130_fd_sc_hd__clkbuf_4 _5576_ (.A(_2631_),
    .X(_2632_));
 sky130_fd_sc_hd__or2_1 _5577_ (.A(_2443_),
    .B(_2334_),
    .X(_2633_));
 sky130_fd_sc_hd__buf_2 _5578_ (.A(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__and3_1 _5579_ (.A(_2473_),
    .B(\dmmu0.page_table[12][0] ),
    .C(_2634_),
    .X(_2635_));
 sky130_fd_sc_hd__a21o_1 _5580_ (.A1(_2211_),
    .A2(_2632_),
    .B1(_2635_),
    .X(_0198_));
 sky130_fd_sc_hd__and3_1 _5581_ (.A(_2473_),
    .B(\dmmu0.page_table[12][1] ),
    .C(_2634_),
    .X(_2636_));
 sky130_fd_sc_hd__a21o_1 _5582_ (.A1(_2224_),
    .A2(_2632_),
    .B1(_2636_),
    .X(_0199_));
 sky130_fd_sc_hd__and3_1 _5583_ (.A(_2473_),
    .B(\dmmu0.page_table[12][2] ),
    .C(_2634_),
    .X(_2637_));
 sky130_fd_sc_hd__a21o_1 _5584_ (.A1(_2227_),
    .A2(_2632_),
    .B1(_2637_),
    .X(_0200_));
 sky130_fd_sc_hd__and3_1 _5585_ (.A(_2473_),
    .B(\dmmu0.page_table[12][3] ),
    .C(_2634_),
    .X(_2638_));
 sky130_fd_sc_hd__a21o_1 _5586_ (.A1(_2230_),
    .A2(_2632_),
    .B1(_2638_),
    .X(_0201_));
 sky130_fd_sc_hd__and3_1 _5587_ (.A(_2473_),
    .B(\dmmu0.page_table[12][4] ),
    .C(_2634_),
    .X(_2639_));
 sky130_fd_sc_hd__a21o_1 _5588_ (.A1(_2233_),
    .A2(_2632_),
    .B1(_2639_),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_4 _5589_ (.A(_2370_),
    .X(_2640_));
 sky130_fd_sc_hd__and3_1 _5590_ (.A(_2640_),
    .B(\dmmu0.page_table[12][5] ),
    .C(_2634_),
    .X(_2641_));
 sky130_fd_sc_hd__a21o_1 _5591_ (.A1(_2236_),
    .A2(_2632_),
    .B1(_2641_),
    .X(_0203_));
 sky130_fd_sc_hd__and3_1 _5592_ (.A(_2640_),
    .B(\dmmu0.page_table[12][6] ),
    .C(_2634_),
    .X(_2642_));
 sky130_fd_sc_hd__a21o_1 _5593_ (.A1(_2240_),
    .A2(_2632_),
    .B1(_2642_),
    .X(_0204_));
 sky130_fd_sc_hd__and3_1 _5594_ (.A(_2640_),
    .B(\dmmu0.page_table[12][7] ),
    .C(_2634_),
    .X(_2643_));
 sky130_fd_sc_hd__a21o_1 _5595_ (.A1(_2243_),
    .A2(_2632_),
    .B1(_2643_),
    .X(_0205_));
 sky130_fd_sc_hd__and3_1 _5596_ (.A(_2640_),
    .B(\dmmu0.page_table[12][8] ),
    .C(_2634_),
    .X(_2644_));
 sky130_fd_sc_hd__a21o_1 _5597_ (.A1(_2245_),
    .A2(_2632_),
    .B1(_2644_),
    .X(_0206_));
 sky130_fd_sc_hd__and3_1 _5598_ (.A(_2640_),
    .B(\dmmu0.page_table[12][9] ),
    .C(_2634_),
    .X(_2645_));
 sky130_fd_sc_hd__a21o_1 _5599_ (.A1(_2247_),
    .A2(_2632_),
    .B1(_2645_),
    .X(_0207_));
 sky130_fd_sc_hd__and3_1 _5600_ (.A(_2640_),
    .B(\dmmu0.page_table[12][10] ),
    .C(_2633_),
    .X(_2646_));
 sky130_fd_sc_hd__a21o_1 _5601_ (.A1(_2249_),
    .A2(_2631_),
    .B1(_2646_),
    .X(_0208_));
 sky130_fd_sc_hd__and3_1 _5602_ (.A(_2640_),
    .B(\dmmu0.page_table[12][11] ),
    .C(_2633_),
    .X(_2647_));
 sky130_fd_sc_hd__a21o_1 _5603_ (.A1(_2251_),
    .A2(_2631_),
    .B1(_2647_),
    .X(_0209_));
 sky130_fd_sc_hd__and3_1 _5604_ (.A(_2640_),
    .B(\dmmu0.page_table[12][12] ),
    .C(_2633_),
    .X(_2648_));
 sky130_fd_sc_hd__a21o_1 _5605_ (.A1(_2253_),
    .A2(_2631_),
    .B1(_2648_),
    .X(_0210_));
 sky130_fd_sc_hd__nor2_1 _5606_ (.A(_2217_),
    .B(_2296_),
    .Y(_2649_));
 sky130_fd_sc_hd__clkbuf_4 _5607_ (.A(_2649_),
    .X(_2650_));
 sky130_fd_sc_hd__or2_1 _5608_ (.A(_2443_),
    .B(_2296_),
    .X(_2651_));
 sky130_fd_sc_hd__buf_2 _5609_ (.A(_2651_),
    .X(_2652_));
 sky130_fd_sc_hd__and3_1 _5610_ (.A(_2640_),
    .B(\dmmu0.page_table[15][0] ),
    .C(_2652_),
    .X(_2653_));
 sky130_fd_sc_hd__a21o_1 _5611_ (.A1(_2211_),
    .A2(_2650_),
    .B1(_2653_),
    .X(_0211_));
 sky130_fd_sc_hd__and3_1 _5612_ (.A(_2640_),
    .B(\dmmu0.page_table[15][1] ),
    .C(_2652_),
    .X(_2654_));
 sky130_fd_sc_hd__a21o_1 _5613_ (.A1(_2224_),
    .A2(_2650_),
    .B1(_2654_),
    .X(_0212_));
 sky130_fd_sc_hd__clkbuf_4 _5614_ (.A(_2370_),
    .X(_2655_));
 sky130_fd_sc_hd__and3_1 _5615_ (.A(_2655_),
    .B(\dmmu0.page_table[15][2] ),
    .C(_2652_),
    .X(_2656_));
 sky130_fd_sc_hd__a21o_1 _5616_ (.A1(_2227_),
    .A2(_2650_),
    .B1(_2656_),
    .X(_0213_));
 sky130_fd_sc_hd__and3_1 _5617_ (.A(_2655_),
    .B(\dmmu0.page_table[15][3] ),
    .C(_2652_),
    .X(_2657_));
 sky130_fd_sc_hd__a21o_1 _5618_ (.A1(_2230_),
    .A2(_2650_),
    .B1(_2657_),
    .X(_0214_));
 sky130_fd_sc_hd__and3_1 _5619_ (.A(_2655_),
    .B(\dmmu0.page_table[15][4] ),
    .C(_2652_),
    .X(_2658_));
 sky130_fd_sc_hd__a21o_1 _5620_ (.A1(_2233_),
    .A2(_2650_),
    .B1(_2658_),
    .X(_0215_));
 sky130_fd_sc_hd__and3_1 _5621_ (.A(_2655_),
    .B(\dmmu0.page_table[15][5] ),
    .C(_2652_),
    .X(_2659_));
 sky130_fd_sc_hd__a21o_1 _5622_ (.A1(_2236_),
    .A2(_2650_),
    .B1(_2659_),
    .X(_0216_));
 sky130_fd_sc_hd__and3_1 _5623_ (.A(_2655_),
    .B(\dmmu0.page_table[15][6] ),
    .C(_2652_),
    .X(_2660_));
 sky130_fd_sc_hd__a21o_1 _5624_ (.A1(_2240_),
    .A2(_2650_),
    .B1(_2660_),
    .X(_0217_));
 sky130_fd_sc_hd__and3_1 _5625_ (.A(_2655_),
    .B(\dmmu0.page_table[15][7] ),
    .C(_2652_),
    .X(_2661_));
 sky130_fd_sc_hd__a21o_1 _5626_ (.A1(_2243_),
    .A2(_2650_),
    .B1(_2661_),
    .X(_0218_));
 sky130_fd_sc_hd__and3_1 _5627_ (.A(_2655_),
    .B(\dmmu0.page_table[15][8] ),
    .C(_2652_),
    .X(_2662_));
 sky130_fd_sc_hd__a21o_1 _5628_ (.A1(_2245_),
    .A2(_2650_),
    .B1(_2662_),
    .X(_0219_));
 sky130_fd_sc_hd__and3_1 _5629_ (.A(_2655_),
    .B(\dmmu0.page_table[15][9] ),
    .C(_2652_),
    .X(_2663_));
 sky130_fd_sc_hd__a21o_1 _5630_ (.A1(_2247_),
    .A2(_2650_),
    .B1(_2663_),
    .X(_0220_));
 sky130_fd_sc_hd__and3_1 _5631_ (.A(_2655_),
    .B(\dmmu0.page_table[15][10] ),
    .C(_2651_),
    .X(_2664_));
 sky130_fd_sc_hd__a21o_1 _5632_ (.A1(_2249_),
    .A2(_2649_),
    .B1(_2664_),
    .X(_0221_));
 sky130_fd_sc_hd__and3_1 _5633_ (.A(_2655_),
    .B(\dmmu0.page_table[15][11] ),
    .C(_2651_),
    .X(_2665_));
 sky130_fd_sc_hd__a21o_1 _5634_ (.A1(_2251_),
    .A2(_2649_),
    .B1(_2665_),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_4 _5635_ (.A(_2370_),
    .X(_2666_));
 sky130_fd_sc_hd__and3_1 _5636_ (.A(_2666_),
    .B(\dmmu0.page_table[15][12] ),
    .C(_2651_),
    .X(_2667_));
 sky130_fd_sc_hd__a21o_1 _5637_ (.A1(_2253_),
    .A2(_2649_),
    .B1(_2667_),
    .X(_0223_));
 sky130_fd_sc_hd__nor2_1 _5638_ (.A(_1914_),
    .B(_2217_),
    .Y(_2668_));
 sky130_fd_sc_hd__buf_4 _5639_ (.A(_2668_),
    .X(_2669_));
 sky130_fd_sc_hd__or2_2 _5640_ (.A(_1914_),
    .B(_2215_),
    .X(_2670_));
 sky130_fd_sc_hd__clkbuf_4 _5641_ (.A(_2670_),
    .X(_2671_));
 sky130_fd_sc_hd__and3_1 _5642_ (.A(_2666_),
    .B(\dmmu0.page_table[11][0] ),
    .C(_2671_),
    .X(_2672_));
 sky130_fd_sc_hd__a21o_1 _5643_ (.A1(_2211_),
    .A2(_2669_),
    .B1(_2672_),
    .X(_0224_));
 sky130_fd_sc_hd__and3_1 _5644_ (.A(_2666_),
    .B(\dmmu0.page_table[11][1] ),
    .C(_2671_),
    .X(_2673_));
 sky130_fd_sc_hd__a21o_1 _5645_ (.A1(_2224_),
    .A2(_2669_),
    .B1(_2673_),
    .X(_0225_));
 sky130_fd_sc_hd__and3_1 _5646_ (.A(_2666_),
    .B(\dmmu0.page_table[11][2] ),
    .C(_2671_),
    .X(_2674_));
 sky130_fd_sc_hd__a21o_1 _5647_ (.A1(_2227_),
    .A2(_2669_),
    .B1(_2674_),
    .X(_0226_));
 sky130_fd_sc_hd__and3_1 _5648_ (.A(_2666_),
    .B(\dmmu0.page_table[11][3] ),
    .C(_2671_),
    .X(_2675_));
 sky130_fd_sc_hd__a21o_1 _5649_ (.A1(_2230_),
    .A2(_2669_),
    .B1(_2675_),
    .X(_0227_));
 sky130_fd_sc_hd__and3_1 _5650_ (.A(_2666_),
    .B(\dmmu0.page_table[11][4] ),
    .C(_2671_),
    .X(_2676_));
 sky130_fd_sc_hd__a21o_1 _5651_ (.A1(_2233_),
    .A2(_2669_),
    .B1(_2676_),
    .X(_0228_));
 sky130_fd_sc_hd__and3_1 _5652_ (.A(_2666_),
    .B(\dmmu0.page_table[11][5] ),
    .C(_2671_),
    .X(_2677_));
 sky130_fd_sc_hd__a21o_1 _5653_ (.A1(_2236_),
    .A2(_2669_),
    .B1(_2677_),
    .X(_0229_));
 sky130_fd_sc_hd__and3_1 _5654_ (.A(_2666_),
    .B(\dmmu0.page_table[11][6] ),
    .C(_2671_),
    .X(_2678_));
 sky130_fd_sc_hd__a21o_1 _5655_ (.A1(_2240_),
    .A2(_2669_),
    .B1(_2678_),
    .X(_0230_));
 sky130_fd_sc_hd__and3_1 _5656_ (.A(_2666_),
    .B(\dmmu0.page_table[11][7] ),
    .C(_2671_),
    .X(_2679_));
 sky130_fd_sc_hd__a21o_1 _5657_ (.A1(_2243_),
    .A2(_2669_),
    .B1(_2679_),
    .X(_0231_));
 sky130_fd_sc_hd__and3_1 _5658_ (.A(_2666_),
    .B(\dmmu0.page_table[11][8] ),
    .C(_2671_),
    .X(_2680_));
 sky130_fd_sc_hd__a21o_1 _5659_ (.A1(_2245_),
    .A2(_2669_),
    .B1(_2680_),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_4 _5660_ (.A(_1896_),
    .X(_2681_));
 sky130_fd_sc_hd__clkbuf_4 _5661_ (.A(_2681_),
    .X(_2682_));
 sky130_fd_sc_hd__and3_1 _5662_ (.A(_2682_),
    .B(\dmmu0.page_table[11][9] ),
    .C(_2671_),
    .X(_2683_));
 sky130_fd_sc_hd__a21o_1 _5663_ (.A1(_2247_),
    .A2(_2669_),
    .B1(_2683_),
    .X(_0233_));
 sky130_fd_sc_hd__and3_1 _5664_ (.A(_2682_),
    .B(\dmmu0.page_table[11][10] ),
    .C(_2670_),
    .X(_2684_));
 sky130_fd_sc_hd__a21o_1 _5665_ (.A1(_2249_),
    .A2(_2668_),
    .B1(_2684_),
    .X(_0234_));
 sky130_fd_sc_hd__and3_1 _5666_ (.A(_2682_),
    .B(\dmmu0.page_table[11][11] ),
    .C(_2670_),
    .X(_2685_));
 sky130_fd_sc_hd__a21o_1 _5667_ (.A1(_2251_),
    .A2(_2668_),
    .B1(_2685_),
    .X(_0235_));
 sky130_fd_sc_hd__and3_1 _5668_ (.A(_2682_),
    .B(\dmmu0.page_table[11][12] ),
    .C(_2670_),
    .X(_2686_));
 sky130_fd_sc_hd__a21o_1 _5669_ (.A1(_2253_),
    .A2(_2668_),
    .B1(_2686_),
    .X(_0236_));
 sky130_fd_sc_hd__clkinv_2 _5670_ (.A(net86),
    .Y(_2687_));
 sky130_fd_sc_hd__or4_2 _5671_ (.A(net710),
    .B(_2687_),
    .C(_1918_),
    .D(_2212_),
    .X(_2688_));
 sky130_fd_sc_hd__or2_1 _5672_ (.A(_1917_),
    .B(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__buf_4 _5673_ (.A(_2689_),
    .X(_2690_));
 sky130_fd_sc_hd__mux2_1 _5674_ (.A0(_2210_),
    .A1(\immu_0.high_addr_off[0] ),
    .S(_2690_),
    .X(_2691_));
 sky130_fd_sc_hd__clkbuf_1 _5675_ (.A(_2691_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _5676_ (.A0(_1928_),
    .A1(\immu_0.high_addr_off[1] ),
    .S(_2690_),
    .X(_2692_));
 sky130_fd_sc_hd__clkbuf_1 _5677_ (.A(_2692_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _5678_ (.A0(_2226_),
    .A1(\immu_0.high_addr_off[2] ),
    .S(_2690_),
    .X(_2693_));
 sky130_fd_sc_hd__clkbuf_1 _5679_ (.A(_2693_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _5680_ (.A0(_2229_),
    .A1(\immu_0.high_addr_off[3] ),
    .S(_2690_),
    .X(_2694_));
 sky130_fd_sc_hd__clkbuf_1 _5681_ (.A(_2694_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _5682_ (.A0(_2232_),
    .A1(\immu_0.high_addr_off[4] ),
    .S(_2690_),
    .X(_2695_));
 sky130_fd_sc_hd__clkbuf_1 _5683_ (.A(_2695_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _5684_ (.A0(_2235_),
    .A1(\immu_0.high_addr_off[5] ),
    .S(_2690_),
    .X(_2696_));
 sky130_fd_sc_hd__clkbuf_1 _5685_ (.A(_2696_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _5686_ (.A0(_2239_),
    .A1(\immu_0.high_addr_off[6] ),
    .S(_2690_),
    .X(_2697_));
 sky130_fd_sc_hd__clkbuf_1 _5687_ (.A(_2697_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5688_ (.A0(_2242_),
    .A1(\immu_0.high_addr_off[7] ),
    .S(_2690_),
    .X(_2698_));
 sky130_fd_sc_hd__clkbuf_1 _5689_ (.A(_2698_),
    .X(_0244_));
 sky130_fd_sc_hd__nor2_1 _5690_ (.A(_2217_),
    .B(_2605_),
    .Y(_2699_));
 sky130_fd_sc_hd__clkbuf_4 _5691_ (.A(_2699_),
    .X(_2700_));
 sky130_fd_sc_hd__or2_1 _5692_ (.A(_2443_),
    .B(_2605_),
    .X(_2701_));
 sky130_fd_sc_hd__buf_2 _5693_ (.A(_2701_),
    .X(_2702_));
 sky130_fd_sc_hd__and3_1 _5694_ (.A(_2682_),
    .B(\dmmu0.page_table[2][0] ),
    .C(_2702_),
    .X(_2703_));
 sky130_fd_sc_hd__a21o_1 _5695_ (.A1(_2211_),
    .A2(_2700_),
    .B1(_2703_),
    .X(_0245_));
 sky130_fd_sc_hd__and3_1 _5696_ (.A(_2682_),
    .B(\dmmu0.page_table[2][1] ),
    .C(_2702_),
    .X(_2704_));
 sky130_fd_sc_hd__a21o_1 _5697_ (.A1(_2224_),
    .A2(_2700_),
    .B1(_2704_),
    .X(_0246_));
 sky130_fd_sc_hd__and3_1 _5698_ (.A(_2682_),
    .B(\dmmu0.page_table[2][2] ),
    .C(_2702_),
    .X(_2705_));
 sky130_fd_sc_hd__a21o_1 _5699_ (.A1(_2227_),
    .A2(_2700_),
    .B1(_2705_),
    .X(_0247_));
 sky130_fd_sc_hd__and3_1 _5700_ (.A(_2682_),
    .B(\dmmu0.page_table[2][3] ),
    .C(_2702_),
    .X(_2706_));
 sky130_fd_sc_hd__a21o_1 _5701_ (.A1(_2230_),
    .A2(_2700_),
    .B1(_2706_),
    .X(_0248_));
 sky130_fd_sc_hd__and3_1 _5702_ (.A(_2682_),
    .B(\dmmu0.page_table[2][4] ),
    .C(_2702_),
    .X(_2707_));
 sky130_fd_sc_hd__a21o_1 _5703_ (.A1(_2233_),
    .A2(_2700_),
    .B1(_2707_),
    .X(_0249_));
 sky130_fd_sc_hd__and3_1 _5704_ (.A(_2682_),
    .B(\dmmu0.page_table[2][5] ),
    .C(_2702_),
    .X(_2708_));
 sky130_fd_sc_hd__a21o_1 _5705_ (.A1(_2236_),
    .A2(_2700_),
    .B1(_2708_),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_4 _5706_ (.A(_2681_),
    .X(_2709_));
 sky130_fd_sc_hd__and3_1 _5707_ (.A(_2709_),
    .B(\dmmu0.page_table[2][6] ),
    .C(_2702_),
    .X(_2710_));
 sky130_fd_sc_hd__a21o_1 _5708_ (.A1(_2240_),
    .A2(_2700_),
    .B1(_2710_),
    .X(_0251_));
 sky130_fd_sc_hd__and3_1 _5709_ (.A(_2709_),
    .B(\dmmu0.page_table[2][7] ),
    .C(_2702_),
    .X(_2711_));
 sky130_fd_sc_hd__a21o_1 _5710_ (.A1(_2243_),
    .A2(_2700_),
    .B1(_2711_),
    .X(_0252_));
 sky130_fd_sc_hd__and3_1 _5711_ (.A(_2709_),
    .B(\dmmu0.page_table[2][8] ),
    .C(_2702_),
    .X(_2712_));
 sky130_fd_sc_hd__a21o_1 _5712_ (.A1(_2245_),
    .A2(_2700_),
    .B1(_2712_),
    .X(_0253_));
 sky130_fd_sc_hd__and3_1 _5713_ (.A(_2709_),
    .B(\dmmu0.page_table[2][9] ),
    .C(_2702_),
    .X(_2713_));
 sky130_fd_sc_hd__a21o_1 _5714_ (.A1(_2247_),
    .A2(_2700_),
    .B1(_2713_),
    .X(_0254_));
 sky130_fd_sc_hd__and3_1 _5715_ (.A(_2709_),
    .B(\dmmu0.page_table[2][10] ),
    .C(_2701_),
    .X(_2714_));
 sky130_fd_sc_hd__a21o_1 _5716_ (.A1(_2249_),
    .A2(_2699_),
    .B1(_2714_),
    .X(_0255_));
 sky130_fd_sc_hd__and3_1 _5717_ (.A(_2709_),
    .B(\dmmu0.page_table[2][11] ),
    .C(_2701_),
    .X(_2715_));
 sky130_fd_sc_hd__a21o_1 _5718_ (.A1(_2251_),
    .A2(_2699_),
    .B1(_2715_),
    .X(_0256_));
 sky130_fd_sc_hd__and3_1 _5719_ (.A(_2709_),
    .B(\dmmu0.page_table[2][12] ),
    .C(_2701_),
    .X(_2716_));
 sky130_fd_sc_hd__a21o_1 _5720_ (.A1(_2253_),
    .A2(_2699_),
    .B1(_2716_),
    .X(_0257_));
 sky130_fd_sc_hd__a21bo_1 _5721_ (.A1(_1579_),
    .A2(net379),
    .B1_N(net325),
    .X(_2717_));
 sky130_fd_sc_hd__o211a_1 _5722_ (.A1(_1579_),
    .A2(net379),
    .B1(_2717_),
    .C1(_1911_),
    .X(_0258_));
 sky130_fd_sc_hd__inv_2 _5723_ (.A(net191),
    .Y(_2718_));
 sky130_fd_sc_hd__or4_4 _5724_ (.A(net710),
    .B(_2718_),
    .C(_1955_),
    .D(_2272_),
    .X(_2719_));
 sky130_fd_sc_hd__nor2_8 _5725_ (.A(_1997_),
    .B(_2719_),
    .Y(_2720_));
 sky130_fd_sc_hd__mux2_1 _5726_ (.A0(\immu_1.high_addr_off[0] ),
    .A1(_1995_),
    .S(_2720_),
    .X(_2721_));
 sky130_fd_sc_hd__clkbuf_1 _5727_ (.A(_2721_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5728_ (.A0(\immu_1.high_addr_off[1] ),
    .A1(_1967_),
    .S(_2720_),
    .X(_2722_));
 sky130_fd_sc_hd__clkbuf_1 _5729_ (.A(_2722_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5730_ (.A0(\immu_1.high_addr_off[2] ),
    .A1(_1972_),
    .S(_2720_),
    .X(_2723_));
 sky130_fd_sc_hd__clkbuf_1 _5731_ (.A(_2723_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5732_ (.A0(\immu_1.high_addr_off[3] ),
    .A1(_1974_),
    .S(_2720_),
    .X(_2724_));
 sky130_fd_sc_hd__clkbuf_1 _5733_ (.A(_2724_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5734_ (.A0(\immu_1.high_addr_off[4] ),
    .A1(_1977_),
    .S(_2720_),
    .X(_2725_));
 sky130_fd_sc_hd__clkbuf_1 _5735_ (.A(_2725_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5736_ (.A0(\immu_1.high_addr_off[5] ),
    .A1(_1979_),
    .S(_2720_),
    .X(_2726_));
 sky130_fd_sc_hd__clkbuf_1 _5737_ (.A(_2726_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _5738_ (.A0(\immu_1.high_addr_off[6] ),
    .A1(_1981_),
    .S(_2720_),
    .X(_2727_));
 sky130_fd_sc_hd__clkbuf_1 _5739_ (.A(_2727_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _5740_ (.A0(\immu_1.high_addr_off[7] ),
    .A1(_1983_),
    .S(_2720_),
    .X(_2728_));
 sky130_fd_sc_hd__clkbuf_1 _5741_ (.A(_2728_),
    .X(_0266_));
 sky130_fd_sc_hd__nor2_2 _5742_ (.A(_2216_),
    .B(_2572_),
    .Y(_2729_));
 sky130_fd_sc_hd__clkbuf_4 _5743_ (.A(_2729_),
    .X(_2730_));
 sky130_fd_sc_hd__or2_1 _5744_ (.A(_2443_),
    .B(_2572_),
    .X(_2731_));
 sky130_fd_sc_hd__buf_2 _5745_ (.A(_2731_),
    .X(_2732_));
 sky130_fd_sc_hd__and3_1 _5746_ (.A(_2709_),
    .B(\dmmu0.page_table[4][0] ),
    .C(_2732_),
    .X(_2733_));
 sky130_fd_sc_hd__a21o_1 _5747_ (.A1(_2210_),
    .A2(_2730_),
    .B1(_2733_),
    .X(_0267_));
 sky130_fd_sc_hd__and3_1 _5748_ (.A(_2709_),
    .B(\dmmu0.page_table[4][1] ),
    .C(_2732_),
    .X(_2734_));
 sky130_fd_sc_hd__a21o_1 _5749_ (.A1(_2223_),
    .A2(_2730_),
    .B1(_2734_),
    .X(_0268_));
 sky130_fd_sc_hd__and3_1 _5750_ (.A(_2709_),
    .B(\dmmu0.page_table[4][2] ),
    .C(_2732_),
    .X(_2735_));
 sky130_fd_sc_hd__a21o_1 _5751_ (.A1(_2226_),
    .A2(_2730_),
    .B1(_2735_),
    .X(_0269_));
 sky130_fd_sc_hd__clkbuf_4 _5752_ (.A(_2681_),
    .X(_2736_));
 sky130_fd_sc_hd__and3_1 _5753_ (.A(_2736_),
    .B(\dmmu0.page_table[4][3] ),
    .C(_2732_),
    .X(_2737_));
 sky130_fd_sc_hd__a21o_1 _5754_ (.A1(_2229_),
    .A2(_2730_),
    .B1(_2737_),
    .X(_0270_));
 sky130_fd_sc_hd__and3_1 _5755_ (.A(_2736_),
    .B(\dmmu0.page_table[4][4] ),
    .C(_2732_),
    .X(_2738_));
 sky130_fd_sc_hd__a21o_1 _5756_ (.A1(_2232_),
    .A2(_2730_),
    .B1(_2738_),
    .X(_0271_));
 sky130_fd_sc_hd__and3_1 _5757_ (.A(_2736_),
    .B(\dmmu0.page_table[4][5] ),
    .C(_2732_),
    .X(_2739_));
 sky130_fd_sc_hd__a21o_1 _5758_ (.A1(_2235_),
    .A2(_2730_),
    .B1(_2739_),
    .X(_0272_));
 sky130_fd_sc_hd__and3_1 _5759_ (.A(_2736_),
    .B(\dmmu0.page_table[4][6] ),
    .C(_2732_),
    .X(_2740_));
 sky130_fd_sc_hd__a21o_1 _5760_ (.A1(_2239_),
    .A2(_2730_),
    .B1(_2740_),
    .X(_0273_));
 sky130_fd_sc_hd__and3_1 _5761_ (.A(_2736_),
    .B(\dmmu0.page_table[4][7] ),
    .C(_2732_),
    .X(_2741_));
 sky130_fd_sc_hd__a21o_1 _5762_ (.A1(_2242_),
    .A2(_2730_),
    .B1(_2741_),
    .X(_0274_));
 sky130_fd_sc_hd__and3_1 _5763_ (.A(_2736_),
    .B(\dmmu0.page_table[4][8] ),
    .C(_2732_),
    .X(_2742_));
 sky130_fd_sc_hd__a21o_1 _5764_ (.A1(_1946_),
    .A2(_2730_),
    .B1(_2742_),
    .X(_0275_));
 sky130_fd_sc_hd__and3_1 _5765_ (.A(_2736_),
    .B(\dmmu0.page_table[4][9] ),
    .C(_2732_),
    .X(_2743_));
 sky130_fd_sc_hd__a21o_1 _5766_ (.A1(_1948_),
    .A2(_2730_),
    .B1(_2743_),
    .X(_0276_));
 sky130_fd_sc_hd__and3_1 _5767_ (.A(_2736_),
    .B(\dmmu0.page_table[4][10] ),
    .C(_2731_),
    .X(_2744_));
 sky130_fd_sc_hd__a21o_1 _5768_ (.A1(_1950_),
    .A2(_2729_),
    .B1(_2744_),
    .X(_0277_));
 sky130_fd_sc_hd__and3_1 _5769_ (.A(_2736_),
    .B(\dmmu0.page_table[4][11] ),
    .C(_2731_),
    .X(_2745_));
 sky130_fd_sc_hd__a21o_1 _5770_ (.A1(net94),
    .A2(_2729_),
    .B1(_2745_),
    .X(_0278_));
 sky130_fd_sc_hd__and3_1 _5771_ (.A(_2736_),
    .B(\dmmu0.page_table[4][12] ),
    .C(_2731_),
    .X(_2746_));
 sky130_fd_sc_hd__a21o_1 _5772_ (.A1(net95),
    .A2(_2729_),
    .B1(_2746_),
    .X(_0279_));
 sky130_fd_sc_hd__nor2_2 _5773_ (.A(_2216_),
    .B(_2351_),
    .Y(_2747_));
 sky130_fd_sc_hd__clkbuf_4 _5774_ (.A(_2747_),
    .X(_2748_));
 sky130_fd_sc_hd__buf_2 _5775_ (.A(_2681_),
    .X(_2749_));
 sky130_fd_sc_hd__or2_2 _5776_ (.A(_2443_),
    .B(_2351_),
    .X(_2750_));
 sky130_fd_sc_hd__buf_2 _5777_ (.A(_2750_),
    .X(_2751_));
 sky130_fd_sc_hd__and3_1 _5778_ (.A(_2749_),
    .B(\dmmu0.page_table[13][0] ),
    .C(_2751_),
    .X(_2752_));
 sky130_fd_sc_hd__a21o_1 _5779_ (.A1(_2210_),
    .A2(_2748_),
    .B1(_2752_),
    .X(_0280_));
 sky130_fd_sc_hd__and3_1 _5780_ (.A(_2749_),
    .B(\dmmu0.page_table[13][1] ),
    .C(_2751_),
    .X(_2753_));
 sky130_fd_sc_hd__a21o_1 _5781_ (.A1(_2223_),
    .A2(_2748_),
    .B1(_2753_),
    .X(_0281_));
 sky130_fd_sc_hd__and3_1 _5782_ (.A(_2749_),
    .B(\dmmu0.page_table[13][2] ),
    .C(_2751_),
    .X(_2754_));
 sky130_fd_sc_hd__a21o_1 _5783_ (.A1(_2226_),
    .A2(_2748_),
    .B1(_2754_),
    .X(_0282_));
 sky130_fd_sc_hd__and3_1 _5784_ (.A(_2749_),
    .B(\dmmu0.page_table[13][3] ),
    .C(_2751_),
    .X(_2755_));
 sky130_fd_sc_hd__a21o_1 _5785_ (.A1(_2229_),
    .A2(_2748_),
    .B1(_2755_),
    .X(_0283_));
 sky130_fd_sc_hd__and3_1 _5786_ (.A(_2749_),
    .B(\dmmu0.page_table[13][4] ),
    .C(_2751_),
    .X(_2756_));
 sky130_fd_sc_hd__a21o_1 _5787_ (.A1(_2232_),
    .A2(_2748_),
    .B1(_2756_),
    .X(_0284_));
 sky130_fd_sc_hd__and3_1 _5788_ (.A(_2749_),
    .B(\dmmu0.page_table[13][5] ),
    .C(_2751_),
    .X(_2757_));
 sky130_fd_sc_hd__a21o_1 _5789_ (.A1(_2235_),
    .A2(_2748_),
    .B1(_2757_),
    .X(_0285_));
 sky130_fd_sc_hd__and3_1 _5790_ (.A(_2749_),
    .B(\dmmu0.page_table[13][6] ),
    .C(_2751_),
    .X(_2758_));
 sky130_fd_sc_hd__a21o_1 _5791_ (.A1(_2239_),
    .A2(_2748_),
    .B1(_2758_),
    .X(_0286_));
 sky130_fd_sc_hd__and3_1 _5792_ (.A(_2749_),
    .B(\dmmu0.page_table[13][7] ),
    .C(_2751_),
    .X(_2759_));
 sky130_fd_sc_hd__a21o_1 _5793_ (.A1(_2242_),
    .A2(_2748_),
    .B1(_2759_),
    .X(_0287_));
 sky130_fd_sc_hd__and3_1 _5794_ (.A(_2749_),
    .B(\dmmu0.page_table[13][8] ),
    .C(_2751_),
    .X(_2760_));
 sky130_fd_sc_hd__a21o_1 _5795_ (.A1(_1946_),
    .A2(_2748_),
    .B1(_2760_),
    .X(_0288_));
 sky130_fd_sc_hd__and3_1 _5796_ (.A(_2749_),
    .B(\dmmu0.page_table[13][9] ),
    .C(_2751_),
    .X(_2761_));
 sky130_fd_sc_hd__a21o_1 _5797_ (.A1(_1948_),
    .A2(_2748_),
    .B1(_2761_),
    .X(_0289_));
 sky130_fd_sc_hd__clkbuf_4 _5798_ (.A(_2681_),
    .X(_2762_));
 sky130_fd_sc_hd__and3_1 _5799_ (.A(_2762_),
    .B(\dmmu0.page_table[13][10] ),
    .C(_2750_),
    .X(_2763_));
 sky130_fd_sc_hd__a21o_1 _5800_ (.A1(_1950_),
    .A2(_2747_),
    .B1(_2763_),
    .X(_0290_));
 sky130_fd_sc_hd__and3_1 _5801_ (.A(_2762_),
    .B(\dmmu0.page_table[13][11] ),
    .C(_2750_),
    .X(_2764_));
 sky130_fd_sc_hd__a21o_1 _5802_ (.A1(net94),
    .A2(_2747_),
    .B1(_2764_),
    .X(_0291_));
 sky130_fd_sc_hd__and3_1 _5803_ (.A(_2762_),
    .B(\dmmu0.page_table[13][12] ),
    .C(_2750_),
    .X(_2765_));
 sky130_fd_sc_hd__a21o_1 _5804_ (.A1(net95),
    .A2(_2747_),
    .B1(_2765_),
    .X(_0292_));
 sky130_fd_sc_hd__nor2_1 _5805_ (.A(_2216_),
    .B(_2589_),
    .Y(_2766_));
 sky130_fd_sc_hd__clkbuf_4 _5806_ (.A(_2766_),
    .X(_2767_));
 sky130_fd_sc_hd__or2_1 _5807_ (.A(_2443_),
    .B(_2589_),
    .X(_2768_));
 sky130_fd_sc_hd__buf_2 _5808_ (.A(_2768_),
    .X(_2769_));
 sky130_fd_sc_hd__and3_1 _5809_ (.A(_2762_),
    .B(\dmmu0.page_table[3][0] ),
    .C(_2769_),
    .X(_2770_));
 sky130_fd_sc_hd__a21o_1 _5810_ (.A1(_2210_),
    .A2(_2767_),
    .B1(_2770_),
    .X(_0293_));
 sky130_fd_sc_hd__and3_1 _5811_ (.A(_2762_),
    .B(\dmmu0.page_table[3][1] ),
    .C(_2769_),
    .X(_2771_));
 sky130_fd_sc_hd__a21o_1 _5812_ (.A1(_2223_),
    .A2(_2767_),
    .B1(_2771_),
    .X(_0294_));
 sky130_fd_sc_hd__and3_1 _5813_ (.A(_2762_),
    .B(\dmmu0.page_table[3][2] ),
    .C(_2769_),
    .X(_2772_));
 sky130_fd_sc_hd__a21o_1 _5814_ (.A1(_2226_),
    .A2(_2767_),
    .B1(_2772_),
    .X(_0295_));
 sky130_fd_sc_hd__and3_1 _5815_ (.A(_2762_),
    .B(\dmmu0.page_table[3][3] ),
    .C(_2769_),
    .X(_2773_));
 sky130_fd_sc_hd__a21o_1 _5816_ (.A1(_2229_),
    .A2(_2767_),
    .B1(_2773_),
    .X(_0296_));
 sky130_fd_sc_hd__and3_1 _5817_ (.A(_2762_),
    .B(\dmmu0.page_table[3][4] ),
    .C(_2769_),
    .X(_2774_));
 sky130_fd_sc_hd__a21o_1 _5818_ (.A1(_2232_),
    .A2(_2767_),
    .B1(_2774_),
    .X(_0297_));
 sky130_fd_sc_hd__and3_1 _5819_ (.A(_2762_),
    .B(\dmmu0.page_table[3][5] ),
    .C(_2769_),
    .X(_2775_));
 sky130_fd_sc_hd__a21o_1 _5820_ (.A1(_2235_),
    .A2(_2767_),
    .B1(_2775_),
    .X(_0298_));
 sky130_fd_sc_hd__and3_1 _5821_ (.A(_2762_),
    .B(\dmmu0.page_table[3][6] ),
    .C(_2769_),
    .X(_2776_));
 sky130_fd_sc_hd__a21o_1 _5822_ (.A1(_2239_),
    .A2(_2767_),
    .B1(_2776_),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_4 _5823_ (.A(_2681_),
    .X(_2777_));
 sky130_fd_sc_hd__and3_1 _5824_ (.A(_2777_),
    .B(\dmmu0.page_table[3][7] ),
    .C(_2769_),
    .X(_2778_));
 sky130_fd_sc_hd__a21o_1 _5825_ (.A1(_2242_),
    .A2(_2767_),
    .B1(_2778_),
    .X(_0300_));
 sky130_fd_sc_hd__and3_1 _5826_ (.A(_2777_),
    .B(\dmmu0.page_table[3][8] ),
    .C(_2769_),
    .X(_2779_));
 sky130_fd_sc_hd__a21o_1 _5827_ (.A1(_1946_),
    .A2(_2767_),
    .B1(_2779_),
    .X(_0301_));
 sky130_fd_sc_hd__and3_1 _5828_ (.A(_2777_),
    .B(\dmmu0.page_table[3][9] ),
    .C(_2769_),
    .X(_2780_));
 sky130_fd_sc_hd__a21o_1 _5829_ (.A1(_1948_),
    .A2(_2767_),
    .B1(_2780_),
    .X(_0302_));
 sky130_fd_sc_hd__and3_1 _5830_ (.A(_2777_),
    .B(\dmmu0.page_table[3][10] ),
    .C(_2768_),
    .X(_2781_));
 sky130_fd_sc_hd__a21o_1 _5831_ (.A1(_1950_),
    .A2(_2766_),
    .B1(_2781_),
    .X(_0303_));
 sky130_fd_sc_hd__and3_1 _5832_ (.A(_2777_),
    .B(\dmmu0.page_table[3][11] ),
    .C(_2768_),
    .X(_2782_));
 sky130_fd_sc_hd__a21o_1 _5833_ (.A1(net94),
    .A2(_2766_),
    .B1(_2782_),
    .X(_0304_));
 sky130_fd_sc_hd__and3_1 _5834_ (.A(_2777_),
    .B(\dmmu0.page_table[3][12] ),
    .C(_2768_),
    .X(_2783_));
 sky130_fd_sc_hd__a21o_1 _5835_ (.A1(net95),
    .A2(_2766_),
    .B1(_2783_),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_4 _5836_ (.A(_1958_),
    .X(_2784_));
 sky130_fd_sc_hd__or2_1 _5837_ (.A(_2784_),
    .B(_2278_),
    .X(_2785_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _5838_ (.A(_2785_),
    .X(_2786_));
 sky130_fd_sc_hd__buf_4 _5839_ (.A(_2786_),
    .X(_2787_));
 sky130_fd_sc_hd__nor2_1 _5840_ (.A(_1968_),
    .B(_2278_),
    .Y(_2788_));
 sky130_fd_sc_hd__clkbuf_4 _5841_ (.A(_2788_),
    .X(_2789_));
 sky130_fd_sc_hd__and2_1 _5842_ (.A(_1995_),
    .B(_2789_),
    .X(_2790_));
 sky130_fd_sc_hd__a31o_1 _5843_ (.A1(_2618_),
    .A2(\dmmu1.page_table[15][0] ),
    .A3(_2787_),
    .B1(_2790_),
    .X(_0306_));
 sky130_fd_sc_hd__buf_2 _5844_ (.A(net201),
    .X(_2791_));
 sky130_fd_sc_hd__and2_1 _5845_ (.A(_2791_),
    .B(_2789_),
    .X(_2792_));
 sky130_fd_sc_hd__a31o_1 _5846_ (.A1(_2618_),
    .A2(\dmmu1.page_table[15][1] ),
    .A3(_2787_),
    .B1(_2792_),
    .X(_0307_));
 sky130_fd_sc_hd__buf_2 _5847_ (.A(net202),
    .X(_2793_));
 sky130_fd_sc_hd__and2_1 _5848_ (.A(_2793_),
    .B(_2789_),
    .X(_2794_));
 sky130_fd_sc_hd__a31o_1 _5849_ (.A1(_2618_),
    .A2(\dmmu1.page_table[15][2] ),
    .A3(_2787_),
    .B1(_2794_),
    .X(_0308_));
 sky130_fd_sc_hd__buf_2 _5850_ (.A(net203),
    .X(_2795_));
 sky130_fd_sc_hd__and2_1 _5851_ (.A(_2795_),
    .B(_2789_),
    .X(_2796_));
 sky130_fd_sc_hd__a31o_1 _5852_ (.A1(_2618_),
    .A2(\dmmu1.page_table[15][3] ),
    .A3(_2787_),
    .B1(_2796_),
    .X(_0309_));
 sky130_fd_sc_hd__buf_2 _5853_ (.A(net204),
    .X(_2797_));
 sky130_fd_sc_hd__and2_1 _5854_ (.A(_2797_),
    .B(_2789_),
    .X(_2798_));
 sky130_fd_sc_hd__a31o_1 _5855_ (.A1(_2618_),
    .A2(\dmmu1.page_table[15][4] ),
    .A3(_2787_),
    .B1(_2798_),
    .X(_0310_));
 sky130_fd_sc_hd__buf_2 _5856_ (.A(net205),
    .X(_2799_));
 sky130_fd_sc_hd__and2_1 _5857_ (.A(_2799_),
    .B(_2789_),
    .X(_2800_));
 sky130_fd_sc_hd__a31o_1 _5858_ (.A1(_2618_),
    .A2(\dmmu1.page_table[15][5] ),
    .A3(_2787_),
    .B1(_2800_),
    .X(_0311_));
 sky130_fd_sc_hd__buf_2 _5859_ (.A(net206),
    .X(_2801_));
 sky130_fd_sc_hd__and2_1 _5860_ (.A(_2801_),
    .B(_2789_),
    .X(_2802_));
 sky130_fd_sc_hd__a31o_1 _5861_ (.A1(_2618_),
    .A2(\dmmu1.page_table[15][6] ),
    .A3(_2787_),
    .B1(_2802_),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_4 _5862_ (.A(net207),
    .X(_2803_));
 sky130_fd_sc_hd__and2_1 _5863_ (.A(_2803_),
    .B(_2789_),
    .X(_2804_));
 sky130_fd_sc_hd__a31o_1 _5864_ (.A1(_2618_),
    .A2(\dmmu1.page_table[15][7] ),
    .A3(_2787_),
    .B1(_2804_),
    .X(_0313_));
 sky130_fd_sc_hd__buf_4 _5865_ (.A(_2561_),
    .X(_2805_));
 sky130_fd_sc_hd__and2_1 _5866_ (.A(_1985_),
    .B(_2789_),
    .X(_2806_));
 sky130_fd_sc_hd__a31o_1 _5867_ (.A1(_2805_),
    .A2(\dmmu1.page_table[15][8] ),
    .A3(_2787_),
    .B1(_2806_),
    .X(_0314_));
 sky130_fd_sc_hd__and2_1 _5868_ (.A(_1987_),
    .B(_2789_),
    .X(_2807_));
 sky130_fd_sc_hd__a31o_1 _5869_ (.A1(_2805_),
    .A2(\dmmu1.page_table[15][9] ),
    .A3(_2787_),
    .B1(_2807_),
    .X(_0315_));
 sky130_fd_sc_hd__and2_1 _5870_ (.A(_1989_),
    .B(_2788_),
    .X(_2808_));
 sky130_fd_sc_hd__a31o_1 _5871_ (.A1(_2805_),
    .A2(\dmmu1.page_table[15][10] ),
    .A3(_2786_),
    .B1(_2808_),
    .X(_0316_));
 sky130_fd_sc_hd__and2_1 _5872_ (.A(_1991_),
    .B(_2788_),
    .X(_2809_));
 sky130_fd_sc_hd__a31o_1 _5873_ (.A1(_2805_),
    .A2(\dmmu1.page_table[15][11] ),
    .A3(_2786_),
    .B1(_2809_),
    .X(_0317_));
 sky130_fd_sc_hd__and2_1 _5874_ (.A(_1993_),
    .B(_2788_),
    .X(_2810_));
 sky130_fd_sc_hd__a31o_1 _5875_ (.A1(_2805_),
    .A2(\dmmu1.page_table[15][12] ),
    .A3(_2786_),
    .B1(_2810_),
    .X(_0318_));
 sky130_fd_sc_hd__nor2_1 _5876_ (.A(_2216_),
    .B(_2539_),
    .Y(_2811_));
 sky130_fd_sc_hd__buf_4 _5877_ (.A(_2811_),
    .X(_2812_));
 sky130_fd_sc_hd__or2_1 _5878_ (.A(_2443_),
    .B(_2539_),
    .X(_2813_));
 sky130_fd_sc_hd__clkbuf_4 _5879_ (.A(_2813_),
    .X(_2814_));
 sky130_fd_sc_hd__and3_1 _5880_ (.A(_2777_),
    .B(\dmmu0.page_table[6][0] ),
    .C(_2814_),
    .X(_2815_));
 sky130_fd_sc_hd__a21o_1 _5881_ (.A1(_2210_),
    .A2(_2812_),
    .B1(_2815_),
    .X(_0319_));
 sky130_fd_sc_hd__and3_1 _5882_ (.A(_2777_),
    .B(\dmmu0.page_table[6][1] ),
    .C(_2814_),
    .X(_2816_));
 sky130_fd_sc_hd__a21o_1 _5883_ (.A1(_2223_),
    .A2(_2812_),
    .B1(_2816_),
    .X(_0320_));
 sky130_fd_sc_hd__and3_1 _5884_ (.A(_2777_),
    .B(\dmmu0.page_table[6][2] ),
    .C(_2814_),
    .X(_2817_));
 sky130_fd_sc_hd__a21o_1 _5885_ (.A1(_2226_),
    .A2(_2812_),
    .B1(_2817_),
    .X(_0321_));
 sky130_fd_sc_hd__and3_1 _5886_ (.A(_2777_),
    .B(\dmmu0.page_table[6][3] ),
    .C(_2814_),
    .X(_2818_));
 sky130_fd_sc_hd__a21o_1 _5887_ (.A1(_2229_),
    .A2(_2812_),
    .B1(_2818_),
    .X(_0322_));
 sky130_fd_sc_hd__buf_2 _5888_ (.A(_2681_),
    .X(_2819_));
 sky130_fd_sc_hd__and3_1 _5889_ (.A(_2819_),
    .B(\dmmu0.page_table[6][4] ),
    .C(_2814_),
    .X(_2820_));
 sky130_fd_sc_hd__a21o_1 _5890_ (.A1(_2232_),
    .A2(_2812_),
    .B1(_2820_),
    .X(_0323_));
 sky130_fd_sc_hd__and3_1 _5891_ (.A(_2819_),
    .B(\dmmu0.page_table[6][5] ),
    .C(_2814_),
    .X(_2821_));
 sky130_fd_sc_hd__a21o_1 _5892_ (.A1(_2235_),
    .A2(_2812_),
    .B1(_2821_),
    .X(_0324_));
 sky130_fd_sc_hd__and3_1 _5893_ (.A(_2819_),
    .B(\dmmu0.page_table[6][6] ),
    .C(_2814_),
    .X(_2822_));
 sky130_fd_sc_hd__a21o_1 _5894_ (.A1(_2239_),
    .A2(_2812_),
    .B1(_2822_),
    .X(_0325_));
 sky130_fd_sc_hd__and3_1 _5895_ (.A(_2819_),
    .B(\dmmu0.page_table[6][7] ),
    .C(_2814_),
    .X(_2823_));
 sky130_fd_sc_hd__a21o_1 _5896_ (.A1(_2242_),
    .A2(_2812_),
    .B1(_2823_),
    .X(_0326_));
 sky130_fd_sc_hd__and3_1 _5897_ (.A(_2819_),
    .B(\dmmu0.page_table[6][8] ),
    .C(_2814_),
    .X(_2824_));
 sky130_fd_sc_hd__a21o_1 _5898_ (.A1(_1946_),
    .A2(_2812_),
    .B1(_2824_),
    .X(_0327_));
 sky130_fd_sc_hd__and3_1 _5899_ (.A(_2819_),
    .B(\dmmu0.page_table[6][9] ),
    .C(_2814_),
    .X(_2825_));
 sky130_fd_sc_hd__a21o_1 _5900_ (.A1(_1948_),
    .A2(_2812_),
    .B1(_2825_),
    .X(_0328_));
 sky130_fd_sc_hd__and3_1 _5901_ (.A(_2819_),
    .B(\dmmu0.page_table[6][10] ),
    .C(_2813_),
    .X(_2826_));
 sky130_fd_sc_hd__a21o_1 _5902_ (.A1(_1950_),
    .A2(_2811_),
    .B1(_2826_),
    .X(_0329_));
 sky130_fd_sc_hd__and3_1 _5903_ (.A(_2819_),
    .B(\dmmu0.page_table[6][11] ),
    .C(_2813_),
    .X(_2827_));
 sky130_fd_sc_hd__a21o_1 _5904_ (.A1(net94),
    .A2(_2811_),
    .B1(_2827_),
    .X(_0330_));
 sky130_fd_sc_hd__and3_1 _5905_ (.A(_2819_),
    .B(\dmmu0.page_table[6][12] ),
    .C(_2813_),
    .X(_2828_));
 sky130_fd_sc_hd__a21o_1 _5906_ (.A1(net95),
    .A2(_2811_),
    .B1(_2828_),
    .X(_0331_));
 sky130_fd_sc_hd__nor2_2 _5907_ (.A(_2216_),
    .B(_2555_),
    .Y(_2829_));
 sky130_fd_sc_hd__buf_4 _5908_ (.A(_2829_),
    .X(_2830_));
 sky130_fd_sc_hd__or2_1 _5909_ (.A(_2443_),
    .B(_2555_),
    .X(_2831_));
 sky130_fd_sc_hd__clkbuf_4 _5910_ (.A(_2831_),
    .X(_2832_));
 sky130_fd_sc_hd__and3_1 _5911_ (.A(_2819_),
    .B(\dmmu0.page_table[5][0] ),
    .C(_2832_),
    .X(_2833_));
 sky130_fd_sc_hd__a21o_1 _5912_ (.A1(_2210_),
    .A2(_2830_),
    .B1(_2833_),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_4 _5913_ (.A(_2681_),
    .X(_2834_));
 sky130_fd_sc_hd__and3_1 _5914_ (.A(_2834_),
    .B(\dmmu0.page_table[5][1] ),
    .C(_2832_),
    .X(_2835_));
 sky130_fd_sc_hd__a21o_1 _5915_ (.A1(_2223_),
    .A2(_2830_),
    .B1(_2835_),
    .X(_0333_));
 sky130_fd_sc_hd__and3_1 _5916_ (.A(_2834_),
    .B(\dmmu0.page_table[5][2] ),
    .C(_2832_),
    .X(_2836_));
 sky130_fd_sc_hd__a21o_1 _5917_ (.A1(_2226_),
    .A2(_2830_),
    .B1(_2836_),
    .X(_0334_));
 sky130_fd_sc_hd__and3_1 _5918_ (.A(_2834_),
    .B(\dmmu0.page_table[5][3] ),
    .C(_2832_),
    .X(_2837_));
 sky130_fd_sc_hd__a21o_1 _5919_ (.A1(_2229_),
    .A2(_2830_),
    .B1(_2837_),
    .X(_0335_));
 sky130_fd_sc_hd__and3_1 _5920_ (.A(_2834_),
    .B(\dmmu0.page_table[5][4] ),
    .C(_2832_),
    .X(_2838_));
 sky130_fd_sc_hd__a21o_1 _5921_ (.A1(_2232_),
    .A2(_2830_),
    .B1(_2838_),
    .X(_0336_));
 sky130_fd_sc_hd__and3_1 _5922_ (.A(_2834_),
    .B(\dmmu0.page_table[5][5] ),
    .C(_2832_),
    .X(_2839_));
 sky130_fd_sc_hd__a21o_1 _5923_ (.A1(_2235_),
    .A2(_2830_),
    .B1(_2839_),
    .X(_0337_));
 sky130_fd_sc_hd__and3_1 _5924_ (.A(_2834_),
    .B(\dmmu0.page_table[5][6] ),
    .C(_2832_),
    .X(_2840_));
 sky130_fd_sc_hd__a21o_1 _5925_ (.A1(_2239_),
    .A2(_2830_),
    .B1(_2840_),
    .X(_0338_));
 sky130_fd_sc_hd__and3_1 _5926_ (.A(_2834_),
    .B(\dmmu0.page_table[5][7] ),
    .C(_2832_),
    .X(_2841_));
 sky130_fd_sc_hd__a21o_1 _5927_ (.A1(_2242_),
    .A2(_2830_),
    .B1(_2841_),
    .X(_0339_));
 sky130_fd_sc_hd__and3_1 _5928_ (.A(_2834_),
    .B(\dmmu0.page_table[5][8] ),
    .C(_2832_),
    .X(_2842_));
 sky130_fd_sc_hd__a21o_1 _5929_ (.A1(_1946_),
    .A2(_2830_),
    .B1(_2842_),
    .X(_0340_));
 sky130_fd_sc_hd__and3_1 _5930_ (.A(_2834_),
    .B(\dmmu0.page_table[5][9] ),
    .C(_2832_),
    .X(_2843_));
 sky130_fd_sc_hd__a21o_1 _5931_ (.A1(_1948_),
    .A2(_2830_),
    .B1(_2843_),
    .X(_0341_));
 sky130_fd_sc_hd__and3_1 _5932_ (.A(_2834_),
    .B(\dmmu0.page_table[5][10] ),
    .C(_2831_),
    .X(_2844_));
 sky130_fd_sc_hd__a21o_1 _5933_ (.A1(_1950_),
    .A2(_2829_),
    .B1(_2844_),
    .X(_0342_));
 sky130_fd_sc_hd__buf_2 _5934_ (.A(_2681_),
    .X(_2845_));
 sky130_fd_sc_hd__and3_1 _5935_ (.A(_2845_),
    .B(\dmmu0.page_table[5][11] ),
    .C(_2831_),
    .X(_2846_));
 sky130_fd_sc_hd__a21o_1 _5936_ (.A1(net94),
    .A2(_2829_),
    .B1(_2846_),
    .X(_0343_));
 sky130_fd_sc_hd__and3_1 _5937_ (.A(_2845_),
    .B(\dmmu0.page_table[5][12] ),
    .C(_2831_),
    .X(_2847_));
 sky130_fd_sc_hd__a21o_1 _5938_ (.A1(net95),
    .A2(_2829_),
    .B1(_2847_),
    .X(_0344_));
 sky130_fd_sc_hd__nor2_4 _5939_ (.A(_2214_),
    .B(_2688_),
    .Y(_2848_));
 sky130_fd_sc_hd__mux2_1 _5940_ (.A0(\dmmu0.long_off_reg[0] ),
    .A1(net92),
    .S(_2848_),
    .X(_2849_));
 sky130_fd_sc_hd__clkbuf_1 _5941_ (.A(_2849_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _5942_ (.A0(\dmmu0.long_off_reg[1] ),
    .A1(_1928_),
    .S(_2848_),
    .X(_2850_));
 sky130_fd_sc_hd__clkbuf_1 _5943_ (.A(_2850_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _5944_ (.A0(\dmmu0.long_off_reg[2] ),
    .A1(_1933_),
    .S(_2848_),
    .X(_2851_));
 sky130_fd_sc_hd__clkbuf_1 _5945_ (.A(_2851_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _5946_ (.A0(\dmmu0.long_off_reg[3] ),
    .A1(_1935_),
    .S(_2848_),
    .X(_2852_));
 sky130_fd_sc_hd__clkbuf_1 _5947_ (.A(_2852_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _5948_ (.A0(\dmmu0.long_off_reg[4] ),
    .A1(_1937_),
    .S(_2848_),
    .X(_2853_));
 sky130_fd_sc_hd__clkbuf_1 _5949_ (.A(_2853_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _5950_ (.A0(\dmmu0.long_off_reg[5] ),
    .A1(_1940_),
    .S(_2848_),
    .X(_2854_));
 sky130_fd_sc_hd__clkbuf_1 _5951_ (.A(_2854_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _5952_ (.A0(\dmmu0.long_off_reg[6] ),
    .A1(_1942_),
    .S(_2848_),
    .X(_2855_));
 sky130_fd_sc_hd__clkbuf_1 _5953_ (.A(_2855_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _5954_ (.A0(\dmmu0.long_off_reg[7] ),
    .A1(_1944_),
    .S(_2848_),
    .X(_2856_));
 sky130_fd_sc_hd__clkbuf_1 _5955_ (.A(_2856_),
    .X(_0352_));
 sky130_fd_sc_hd__or2_1 _5956_ (.A(_2784_),
    .B(_2028_),
    .X(_2857_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _5957_ (.A(_2857_),
    .X(_2858_));
 sky130_fd_sc_hd__buf_4 _5958_ (.A(_2858_),
    .X(_2859_));
 sky130_fd_sc_hd__nor2_1 _5959_ (.A(_1968_),
    .B(_2028_),
    .Y(_2860_));
 sky130_fd_sc_hd__clkbuf_4 _5960_ (.A(_2860_),
    .X(_2861_));
 sky130_fd_sc_hd__and2_1 _5961_ (.A(_1995_),
    .B(_2861_),
    .X(_2862_));
 sky130_fd_sc_hd__a31o_1 _5962_ (.A1(_2805_),
    .A2(\dmmu1.page_table[13][0] ),
    .A3(_2859_),
    .B1(_2862_),
    .X(_0353_));
 sky130_fd_sc_hd__and2_1 _5963_ (.A(_2791_),
    .B(_2861_),
    .X(_2863_));
 sky130_fd_sc_hd__a31o_1 _5964_ (.A1(_2805_),
    .A2(\dmmu1.page_table[13][1] ),
    .A3(_2859_),
    .B1(_2863_),
    .X(_0354_));
 sky130_fd_sc_hd__and2_1 _5965_ (.A(_2793_),
    .B(_2861_),
    .X(_2864_));
 sky130_fd_sc_hd__a31o_1 _5966_ (.A1(_2805_),
    .A2(\dmmu1.page_table[13][2] ),
    .A3(_2859_),
    .B1(_2864_),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _5967_ (.A(_2795_),
    .B(_2861_),
    .X(_2865_));
 sky130_fd_sc_hd__a31o_1 _5968_ (.A1(_2805_),
    .A2(\dmmu1.page_table[13][3] ),
    .A3(_2859_),
    .B1(_2865_),
    .X(_0356_));
 sky130_fd_sc_hd__and2_1 _5969_ (.A(_2797_),
    .B(_2861_),
    .X(_2866_));
 sky130_fd_sc_hd__a31o_1 _5970_ (.A1(_2805_),
    .A2(\dmmu1.page_table[13][4] ),
    .A3(_2859_),
    .B1(_2866_),
    .X(_0357_));
 sky130_fd_sc_hd__buf_4 _5971_ (.A(_2561_),
    .X(_2867_));
 sky130_fd_sc_hd__and2_1 _5972_ (.A(_2799_),
    .B(_2861_),
    .X(_2868_));
 sky130_fd_sc_hd__a31o_1 _5973_ (.A1(_2867_),
    .A2(\dmmu1.page_table[13][5] ),
    .A3(_2859_),
    .B1(_2868_),
    .X(_0358_));
 sky130_fd_sc_hd__and2_1 _5974_ (.A(_2801_),
    .B(_2861_),
    .X(_2869_));
 sky130_fd_sc_hd__a31o_1 _5975_ (.A1(_2867_),
    .A2(\dmmu1.page_table[13][6] ),
    .A3(_2859_),
    .B1(_2869_),
    .X(_0359_));
 sky130_fd_sc_hd__and2_1 _5976_ (.A(_2803_),
    .B(_2861_),
    .X(_2870_));
 sky130_fd_sc_hd__a31o_1 _5977_ (.A1(_2867_),
    .A2(\dmmu1.page_table[13][7] ),
    .A3(_2859_),
    .B1(_2870_),
    .X(_0360_));
 sky130_fd_sc_hd__and2_1 _5978_ (.A(_1985_),
    .B(_2861_),
    .X(_2871_));
 sky130_fd_sc_hd__a31o_1 _5979_ (.A1(_2867_),
    .A2(\dmmu1.page_table[13][8] ),
    .A3(_2859_),
    .B1(_2871_),
    .X(_0361_));
 sky130_fd_sc_hd__and2_1 _5980_ (.A(_1987_),
    .B(_2861_),
    .X(_2872_));
 sky130_fd_sc_hd__a31o_1 _5981_ (.A1(_2867_),
    .A2(\dmmu1.page_table[13][9] ),
    .A3(_2859_),
    .B1(_2872_),
    .X(_0362_));
 sky130_fd_sc_hd__and2_1 _5982_ (.A(_1989_),
    .B(_2860_),
    .X(_2873_));
 sky130_fd_sc_hd__a31o_1 _5983_ (.A1(_2867_),
    .A2(\dmmu1.page_table[13][10] ),
    .A3(_2858_),
    .B1(_2873_),
    .X(_0363_));
 sky130_fd_sc_hd__and2_1 _5984_ (.A(_1991_),
    .B(_2860_),
    .X(_2874_));
 sky130_fd_sc_hd__a31o_1 _5985_ (.A1(_2867_),
    .A2(\dmmu1.page_table[13][11] ),
    .A3(_2858_),
    .B1(_2874_),
    .X(_0364_));
 sky130_fd_sc_hd__and2_1 _5986_ (.A(_1993_),
    .B(_2860_),
    .X(_2875_));
 sky130_fd_sc_hd__a31o_1 _5987_ (.A1(_2867_),
    .A2(\dmmu1.page_table[13][12] ),
    .A3(_2858_),
    .B1(_2875_),
    .X(_0365_));
 sky130_fd_sc_hd__or2_1 _5988_ (.A(_2784_),
    .B(_2045_),
    .X(_2876_));
 sky130_fd_sc_hd__clkbuf_2 _5989_ (.A(_2876_),
    .X(_2877_));
 sky130_fd_sc_hd__clkbuf_4 _5990_ (.A(_2877_),
    .X(_2878_));
 sky130_fd_sc_hd__buf_2 _5991_ (.A(net197),
    .X(_2879_));
 sky130_fd_sc_hd__nor2_2 _5992_ (.A(_1968_),
    .B(_2045_),
    .Y(_2880_));
 sky130_fd_sc_hd__buf_2 _5993_ (.A(_2880_),
    .X(_2881_));
 sky130_fd_sc_hd__and2_1 _5994_ (.A(_2879_),
    .B(_2881_),
    .X(_2882_));
 sky130_fd_sc_hd__a31o_1 _5995_ (.A1(_2867_),
    .A2(\dmmu1.page_table[12][0] ),
    .A3(_2878_),
    .B1(_2882_),
    .X(_0366_));
 sky130_fd_sc_hd__and2_1 _5996_ (.A(_2791_),
    .B(_2881_),
    .X(_2883_));
 sky130_fd_sc_hd__a31o_1 _5997_ (.A1(_2867_),
    .A2(\dmmu1.page_table[12][1] ),
    .A3(_2878_),
    .B1(_2883_),
    .X(_0367_));
 sky130_fd_sc_hd__buf_4 _5998_ (.A(_2561_),
    .X(_2884_));
 sky130_fd_sc_hd__and2_1 _5999_ (.A(_2793_),
    .B(_2881_),
    .X(_2885_));
 sky130_fd_sc_hd__a31o_1 _6000_ (.A1(_2884_),
    .A2(\dmmu1.page_table[12][2] ),
    .A3(_2878_),
    .B1(_2885_),
    .X(_0368_));
 sky130_fd_sc_hd__and2_1 _6001_ (.A(_2795_),
    .B(_2881_),
    .X(_2886_));
 sky130_fd_sc_hd__a31o_1 _6002_ (.A1(_2884_),
    .A2(\dmmu1.page_table[12][3] ),
    .A3(_2878_),
    .B1(_2886_),
    .X(_0369_));
 sky130_fd_sc_hd__and2_1 _6003_ (.A(_2797_),
    .B(_2881_),
    .X(_2887_));
 sky130_fd_sc_hd__a31o_1 _6004_ (.A1(_2884_),
    .A2(\dmmu1.page_table[12][4] ),
    .A3(_2878_),
    .B1(_2887_),
    .X(_0370_));
 sky130_fd_sc_hd__and2_1 _6005_ (.A(_2799_),
    .B(_2881_),
    .X(_2888_));
 sky130_fd_sc_hd__a31o_1 _6006_ (.A1(_2884_),
    .A2(\dmmu1.page_table[12][5] ),
    .A3(_2878_),
    .B1(_2888_),
    .X(_0371_));
 sky130_fd_sc_hd__and2_1 _6007_ (.A(_2801_),
    .B(_2881_),
    .X(_2889_));
 sky130_fd_sc_hd__a31o_1 _6008_ (.A1(_2884_),
    .A2(\dmmu1.page_table[12][6] ),
    .A3(_2878_),
    .B1(_2889_),
    .X(_0372_));
 sky130_fd_sc_hd__and2_1 _6009_ (.A(_2803_),
    .B(_2881_),
    .X(_2890_));
 sky130_fd_sc_hd__a31o_1 _6010_ (.A1(_2884_),
    .A2(\dmmu1.page_table[12][7] ),
    .A3(_2878_),
    .B1(_2890_),
    .X(_0373_));
 sky130_fd_sc_hd__buf_2 _6011_ (.A(net208),
    .X(_2891_));
 sky130_fd_sc_hd__and2_1 _6012_ (.A(_2891_),
    .B(_2881_),
    .X(_2892_));
 sky130_fd_sc_hd__a31o_1 _6013_ (.A1(_2884_),
    .A2(\dmmu1.page_table[12][8] ),
    .A3(_2878_),
    .B1(_2892_),
    .X(_0374_));
 sky130_fd_sc_hd__buf_2 _6014_ (.A(net209),
    .X(_2893_));
 sky130_fd_sc_hd__and2_1 _6015_ (.A(_2893_),
    .B(_2881_),
    .X(_2894_));
 sky130_fd_sc_hd__a31o_1 _6016_ (.A1(_2884_),
    .A2(\dmmu1.page_table[12][9] ),
    .A3(_2878_),
    .B1(_2894_),
    .X(_0375_));
 sky130_fd_sc_hd__buf_2 _6017_ (.A(net198),
    .X(_2895_));
 sky130_fd_sc_hd__and2_1 _6018_ (.A(_2895_),
    .B(_2880_),
    .X(_2896_));
 sky130_fd_sc_hd__a31o_1 _6019_ (.A1(_2884_),
    .A2(\dmmu1.page_table[12][10] ),
    .A3(_2877_),
    .B1(_2896_),
    .X(_0376_));
 sky130_fd_sc_hd__and2_1 _6020_ (.A(_1991_),
    .B(_2880_),
    .X(_2897_));
 sky130_fd_sc_hd__a31o_1 _6021_ (.A1(_2884_),
    .A2(\dmmu1.page_table[12][11] ),
    .A3(_2877_),
    .B1(_2897_),
    .X(_0377_));
 sky130_fd_sc_hd__buf_4 _6022_ (.A(_2561_),
    .X(_2898_));
 sky130_fd_sc_hd__and2_1 _6023_ (.A(_1993_),
    .B(_2880_),
    .X(_2899_));
 sky130_fd_sc_hd__a31o_1 _6024_ (.A1(_2898_),
    .A2(\dmmu1.page_table[12][12] ),
    .A3(_2877_),
    .B1(_2899_),
    .X(_0378_));
 sky130_fd_sc_hd__or2_1 _6025_ (.A(_2784_),
    .B(_2064_),
    .X(_2900_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _6026_ (.A(_2900_),
    .X(_2901_));
 sky130_fd_sc_hd__buf_4 _6027_ (.A(_2901_),
    .X(_2902_));
 sky130_fd_sc_hd__nor2_1 _6028_ (.A(_1968_),
    .B(_2064_),
    .Y(_2903_));
 sky130_fd_sc_hd__clkbuf_4 _6029_ (.A(_2903_),
    .X(_2904_));
 sky130_fd_sc_hd__and2_1 _6030_ (.A(_2879_),
    .B(_2904_),
    .X(_2905_));
 sky130_fd_sc_hd__a31o_1 _6031_ (.A1(_2898_),
    .A2(\dmmu1.page_table[11][0] ),
    .A3(_2902_),
    .B1(_2905_),
    .X(_0379_));
 sky130_fd_sc_hd__and2_1 _6032_ (.A(_2791_),
    .B(_2904_),
    .X(_2906_));
 sky130_fd_sc_hd__a31o_1 _6033_ (.A1(_2898_),
    .A2(\dmmu1.page_table[11][1] ),
    .A3(_2902_),
    .B1(_2906_),
    .X(_0380_));
 sky130_fd_sc_hd__and2_1 _6034_ (.A(_2793_),
    .B(_2904_),
    .X(_2907_));
 sky130_fd_sc_hd__a31o_1 _6035_ (.A1(_2898_),
    .A2(\dmmu1.page_table[11][2] ),
    .A3(_2902_),
    .B1(_2907_),
    .X(_0381_));
 sky130_fd_sc_hd__and2_1 _6036_ (.A(_2795_),
    .B(_2904_),
    .X(_2908_));
 sky130_fd_sc_hd__a31o_1 _6037_ (.A1(_2898_),
    .A2(\dmmu1.page_table[11][3] ),
    .A3(_2902_),
    .B1(_2908_),
    .X(_0382_));
 sky130_fd_sc_hd__and2_1 _6038_ (.A(_2797_),
    .B(_2904_),
    .X(_2909_));
 sky130_fd_sc_hd__a31o_1 _6039_ (.A1(_2898_),
    .A2(\dmmu1.page_table[11][4] ),
    .A3(_2902_),
    .B1(_2909_),
    .X(_0383_));
 sky130_fd_sc_hd__and2_1 _6040_ (.A(_2799_),
    .B(_2904_),
    .X(_2910_));
 sky130_fd_sc_hd__a31o_1 _6041_ (.A1(_2898_),
    .A2(\dmmu1.page_table[11][5] ),
    .A3(_2902_),
    .B1(_2910_),
    .X(_0384_));
 sky130_fd_sc_hd__and2_1 _6042_ (.A(_2801_),
    .B(_2904_),
    .X(_2911_));
 sky130_fd_sc_hd__a31o_1 _6043_ (.A1(_2898_),
    .A2(\dmmu1.page_table[11][6] ),
    .A3(_2902_),
    .B1(_2911_),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _6044_ (.A(_2803_),
    .B(_2904_),
    .X(_2912_));
 sky130_fd_sc_hd__a31o_1 _6045_ (.A1(_2898_),
    .A2(\dmmu1.page_table[11][7] ),
    .A3(_2902_),
    .B1(_2912_),
    .X(_0386_));
 sky130_fd_sc_hd__and2_1 _6046_ (.A(_2891_),
    .B(_2904_),
    .X(_2913_));
 sky130_fd_sc_hd__a31o_1 _6047_ (.A1(_2898_),
    .A2(\dmmu1.page_table[11][8] ),
    .A3(_2902_),
    .B1(_2913_),
    .X(_0387_));
 sky130_fd_sc_hd__buf_4 _6048_ (.A(_2561_),
    .X(_2914_));
 sky130_fd_sc_hd__and2_1 _6049_ (.A(_2893_),
    .B(_2904_),
    .X(_2915_));
 sky130_fd_sc_hd__a31o_1 _6050_ (.A1(_2914_),
    .A2(\dmmu1.page_table[11][9] ),
    .A3(_2902_),
    .B1(_2915_),
    .X(_0388_));
 sky130_fd_sc_hd__and2_1 _6051_ (.A(_2895_),
    .B(_2903_),
    .X(_2916_));
 sky130_fd_sc_hd__a31o_1 _6052_ (.A1(_2914_),
    .A2(\dmmu1.page_table[11][10] ),
    .A3(_2901_),
    .B1(_2916_),
    .X(_0389_));
 sky130_fd_sc_hd__and2_1 _6053_ (.A(_1991_),
    .B(_2903_),
    .X(_2917_));
 sky130_fd_sc_hd__a31o_1 _6054_ (.A1(_2914_),
    .A2(\dmmu1.page_table[11][11] ),
    .A3(_2901_),
    .B1(_2917_),
    .X(_0390_));
 sky130_fd_sc_hd__and2_1 _6055_ (.A(_1993_),
    .B(_2903_),
    .X(_2918_));
 sky130_fd_sc_hd__a31o_1 _6056_ (.A1(_2914_),
    .A2(\dmmu1.page_table[11][12] ),
    .A3(_2901_),
    .B1(_2918_),
    .X(_0391_));
 sky130_fd_sc_hd__buf_2 _6057_ (.A(_1958_),
    .X(_2919_));
 sky130_fd_sc_hd__or2_1 _6058_ (.A(_2919_),
    .B(_2081_),
    .X(_2920_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _6059_ (.A(_2920_),
    .X(_2921_));
 sky130_fd_sc_hd__buf_4 _6060_ (.A(_2921_),
    .X(_2922_));
 sky130_fd_sc_hd__nor2_1 _6061_ (.A(_1968_),
    .B(_2081_),
    .Y(_2923_));
 sky130_fd_sc_hd__clkbuf_4 _6062_ (.A(_2923_),
    .X(_2924_));
 sky130_fd_sc_hd__and2_1 _6063_ (.A(_2879_),
    .B(_2924_),
    .X(_2925_));
 sky130_fd_sc_hd__a31o_1 _6064_ (.A1(_2914_),
    .A2(\dmmu1.page_table[10][0] ),
    .A3(_2922_),
    .B1(_2925_),
    .X(_0392_));
 sky130_fd_sc_hd__and2_1 _6065_ (.A(_2791_),
    .B(_2924_),
    .X(_2926_));
 sky130_fd_sc_hd__a31o_1 _6066_ (.A1(_2914_),
    .A2(\dmmu1.page_table[10][1] ),
    .A3(_2922_),
    .B1(_2926_),
    .X(_0393_));
 sky130_fd_sc_hd__and2_1 _6067_ (.A(_2793_),
    .B(_2924_),
    .X(_2927_));
 sky130_fd_sc_hd__a31o_1 _6068_ (.A1(_2914_),
    .A2(\dmmu1.page_table[10][2] ),
    .A3(_2922_),
    .B1(_2927_),
    .X(_0394_));
 sky130_fd_sc_hd__and2_1 _6069_ (.A(_2795_),
    .B(_2924_),
    .X(_2928_));
 sky130_fd_sc_hd__a31o_1 _6070_ (.A1(_2914_),
    .A2(\dmmu1.page_table[10][3] ),
    .A3(_2922_),
    .B1(_2928_),
    .X(_0395_));
 sky130_fd_sc_hd__and2_1 _6071_ (.A(_2797_),
    .B(_2924_),
    .X(_2929_));
 sky130_fd_sc_hd__a31o_1 _6072_ (.A1(_2914_),
    .A2(\dmmu1.page_table[10][4] ),
    .A3(_2922_),
    .B1(_2929_),
    .X(_0396_));
 sky130_fd_sc_hd__and2_1 _6073_ (.A(_2799_),
    .B(_2924_),
    .X(_2930_));
 sky130_fd_sc_hd__a31o_1 _6074_ (.A1(_2914_),
    .A2(\dmmu1.page_table[10][5] ),
    .A3(_2922_),
    .B1(_2930_),
    .X(_0397_));
 sky130_fd_sc_hd__buf_2 _6075_ (.A(_1897_),
    .X(_2931_));
 sky130_fd_sc_hd__buf_4 _6076_ (.A(_2931_),
    .X(_2932_));
 sky130_fd_sc_hd__and2_1 _6077_ (.A(_2801_),
    .B(_2924_),
    .X(_2933_));
 sky130_fd_sc_hd__a31o_1 _6078_ (.A1(_2932_),
    .A2(\dmmu1.page_table[10][6] ),
    .A3(_2922_),
    .B1(_2933_),
    .X(_0398_));
 sky130_fd_sc_hd__and2_1 _6079_ (.A(_2803_),
    .B(_2924_),
    .X(_2934_));
 sky130_fd_sc_hd__a31o_1 _6080_ (.A1(_2932_),
    .A2(\dmmu1.page_table[10][7] ),
    .A3(_2922_),
    .B1(_2934_),
    .X(_0399_));
 sky130_fd_sc_hd__and2_1 _6081_ (.A(_2891_),
    .B(_2924_),
    .X(_2935_));
 sky130_fd_sc_hd__a31o_1 _6082_ (.A1(_2932_),
    .A2(\dmmu1.page_table[10][8] ),
    .A3(_2922_),
    .B1(_2935_),
    .X(_0400_));
 sky130_fd_sc_hd__and2_1 _6083_ (.A(_2893_),
    .B(_2924_),
    .X(_2936_));
 sky130_fd_sc_hd__a31o_1 _6084_ (.A1(_2932_),
    .A2(\dmmu1.page_table[10][9] ),
    .A3(_2922_),
    .B1(_2936_),
    .X(_0401_));
 sky130_fd_sc_hd__and2_1 _6085_ (.A(_2895_),
    .B(_2923_),
    .X(_2937_));
 sky130_fd_sc_hd__a31o_1 _6086_ (.A1(_2932_),
    .A2(\dmmu1.page_table[10][10] ),
    .A3(_2921_),
    .B1(_2937_),
    .X(_0402_));
 sky130_fd_sc_hd__and2_1 _6087_ (.A(_1991_),
    .B(_2923_),
    .X(_2938_));
 sky130_fd_sc_hd__a31o_1 _6088_ (.A1(_2932_),
    .A2(\dmmu1.page_table[10][11] ),
    .A3(_2921_),
    .B1(_2938_),
    .X(_0403_));
 sky130_fd_sc_hd__and2_1 _6089_ (.A(_1993_),
    .B(_2923_),
    .X(_2939_));
 sky130_fd_sc_hd__a31o_1 _6090_ (.A1(_2932_),
    .A2(\dmmu1.page_table[10][12] ),
    .A3(_2921_),
    .B1(_2939_),
    .X(_0404_));
 sky130_fd_sc_hd__or2_1 _6091_ (.A(_2919_),
    .B(_2099_),
    .X(_2940_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _6092_ (.A(_2940_),
    .X(_2941_));
 sky130_fd_sc_hd__clkbuf_4 _6093_ (.A(_2941_),
    .X(_2942_));
 sky130_fd_sc_hd__nor2_1 _6094_ (.A(_1968_),
    .B(_2099_),
    .Y(_2943_));
 sky130_fd_sc_hd__clkbuf_4 _6095_ (.A(_2943_),
    .X(_2944_));
 sky130_fd_sc_hd__and2_1 _6096_ (.A(_2879_),
    .B(_2944_),
    .X(_2945_));
 sky130_fd_sc_hd__a31o_1 _6097_ (.A1(_2932_),
    .A2(\dmmu1.page_table[9][0] ),
    .A3(_2942_),
    .B1(_2945_),
    .X(_0405_));
 sky130_fd_sc_hd__and2_1 _6098_ (.A(_2791_),
    .B(_2944_),
    .X(_2946_));
 sky130_fd_sc_hd__a31o_1 _6099_ (.A1(_2932_),
    .A2(\dmmu1.page_table[9][1] ),
    .A3(_2942_),
    .B1(_2946_),
    .X(_0406_));
 sky130_fd_sc_hd__and2_1 _6100_ (.A(_2793_),
    .B(_2944_),
    .X(_2947_));
 sky130_fd_sc_hd__a31o_1 _6101_ (.A1(_2932_),
    .A2(\dmmu1.page_table[9][2] ),
    .A3(_2942_),
    .B1(_2947_),
    .X(_0407_));
 sky130_fd_sc_hd__buf_4 _6102_ (.A(_2931_),
    .X(_2948_));
 sky130_fd_sc_hd__and2_1 _6103_ (.A(_2795_),
    .B(_2944_),
    .X(_2949_));
 sky130_fd_sc_hd__a31o_1 _6104_ (.A1(_2948_),
    .A2(\dmmu1.page_table[9][3] ),
    .A3(_2942_),
    .B1(_2949_),
    .X(_0408_));
 sky130_fd_sc_hd__and2_1 _6105_ (.A(_2797_),
    .B(_2944_),
    .X(_2950_));
 sky130_fd_sc_hd__a31o_1 _6106_ (.A1(_2948_),
    .A2(\dmmu1.page_table[9][4] ),
    .A3(_2942_),
    .B1(_2950_),
    .X(_0409_));
 sky130_fd_sc_hd__and2_1 _6107_ (.A(_2799_),
    .B(_2944_),
    .X(_2951_));
 sky130_fd_sc_hd__a31o_1 _6108_ (.A1(_2948_),
    .A2(\dmmu1.page_table[9][5] ),
    .A3(_2942_),
    .B1(_2951_),
    .X(_0410_));
 sky130_fd_sc_hd__and2_1 _6109_ (.A(_2801_),
    .B(_2944_),
    .X(_2952_));
 sky130_fd_sc_hd__a31o_1 _6110_ (.A1(_2948_),
    .A2(\dmmu1.page_table[9][6] ),
    .A3(_2942_),
    .B1(_2952_),
    .X(_0411_));
 sky130_fd_sc_hd__and2_1 _6111_ (.A(_2803_),
    .B(_2944_),
    .X(_2953_));
 sky130_fd_sc_hd__a31o_1 _6112_ (.A1(_2948_),
    .A2(\dmmu1.page_table[9][7] ),
    .A3(_2942_),
    .B1(_2953_),
    .X(_0412_));
 sky130_fd_sc_hd__and2_1 _6113_ (.A(_2891_),
    .B(_2944_),
    .X(_2954_));
 sky130_fd_sc_hd__a31o_1 _6114_ (.A1(_2948_),
    .A2(\dmmu1.page_table[9][8] ),
    .A3(_2942_),
    .B1(_2954_),
    .X(_0413_));
 sky130_fd_sc_hd__and2_1 _6115_ (.A(_2893_),
    .B(_2944_),
    .X(_2955_));
 sky130_fd_sc_hd__a31o_1 _6116_ (.A1(_2948_),
    .A2(\dmmu1.page_table[9][9] ),
    .A3(_2942_),
    .B1(_2955_),
    .X(_0414_));
 sky130_fd_sc_hd__and2_1 _6117_ (.A(_2895_),
    .B(_2943_),
    .X(_2956_));
 sky130_fd_sc_hd__a31o_1 _6118_ (.A1(_2948_),
    .A2(\dmmu1.page_table[9][10] ),
    .A3(_2941_),
    .B1(_2956_),
    .X(_0415_));
 sky130_fd_sc_hd__and2_1 _6119_ (.A(_1991_),
    .B(_2943_),
    .X(_2957_));
 sky130_fd_sc_hd__a31o_1 _6120_ (.A1(_2948_),
    .A2(\dmmu1.page_table[9][11] ),
    .A3(_2941_),
    .B1(_2957_),
    .X(_0416_));
 sky130_fd_sc_hd__and2_1 _6121_ (.A(_1993_),
    .B(_2943_),
    .X(_2958_));
 sky130_fd_sc_hd__a31o_1 _6122_ (.A1(_2948_),
    .A2(\dmmu1.page_table[9][12] ),
    .A3(_2941_),
    .B1(_2958_),
    .X(_0417_));
 sky130_fd_sc_hd__nor2_1 _6123_ (.A(_2216_),
    .B(_2621_),
    .Y(_2959_));
 sky130_fd_sc_hd__clkbuf_4 _6124_ (.A(_2959_),
    .X(_2960_));
 sky130_fd_sc_hd__or2_1 _6125_ (.A(_2215_),
    .B(_2621_),
    .X(_2961_));
 sky130_fd_sc_hd__clkbuf_4 _6126_ (.A(_2961_),
    .X(_2962_));
 sky130_fd_sc_hd__and3_1 _6127_ (.A(_2845_),
    .B(\dmmu0.page_table[1][0] ),
    .C(_2962_),
    .X(_2963_));
 sky130_fd_sc_hd__a21o_1 _6128_ (.A1(_2210_),
    .A2(_2960_),
    .B1(_2963_),
    .X(_0418_));
 sky130_fd_sc_hd__and3_1 _6129_ (.A(_2845_),
    .B(\dmmu0.page_table[1][1] ),
    .C(_2962_),
    .X(_2964_));
 sky130_fd_sc_hd__a21o_1 _6130_ (.A1(_2223_),
    .A2(_2960_),
    .B1(_2964_),
    .X(_0419_));
 sky130_fd_sc_hd__and3_1 _6131_ (.A(_2845_),
    .B(\dmmu0.page_table[1][2] ),
    .C(_2962_),
    .X(_2965_));
 sky130_fd_sc_hd__a21o_1 _6132_ (.A1(_2226_),
    .A2(_2960_),
    .B1(_2965_),
    .X(_0420_));
 sky130_fd_sc_hd__and3_1 _6133_ (.A(_2845_),
    .B(\dmmu0.page_table[1][3] ),
    .C(_2962_),
    .X(_2966_));
 sky130_fd_sc_hd__a21o_1 _6134_ (.A1(_2229_),
    .A2(_2960_),
    .B1(_2966_),
    .X(_0421_));
 sky130_fd_sc_hd__and3_1 _6135_ (.A(_2845_),
    .B(\dmmu0.page_table[1][4] ),
    .C(_2962_),
    .X(_2967_));
 sky130_fd_sc_hd__a21o_1 _6136_ (.A1(_2232_),
    .A2(_2960_),
    .B1(_2967_),
    .X(_0422_));
 sky130_fd_sc_hd__and3_1 _6137_ (.A(_2845_),
    .B(\dmmu0.page_table[1][5] ),
    .C(_2962_),
    .X(_2968_));
 sky130_fd_sc_hd__a21o_1 _6138_ (.A1(_2235_),
    .A2(_2960_),
    .B1(_2968_),
    .X(_0423_));
 sky130_fd_sc_hd__and3_1 _6139_ (.A(_2845_),
    .B(\dmmu0.page_table[1][6] ),
    .C(_2962_),
    .X(_2969_));
 sky130_fd_sc_hd__a21o_1 _6140_ (.A1(_2239_),
    .A2(_2960_),
    .B1(_2969_),
    .X(_0424_));
 sky130_fd_sc_hd__and3_1 _6141_ (.A(_2845_),
    .B(\dmmu0.page_table[1][7] ),
    .C(_2962_),
    .X(_2970_));
 sky130_fd_sc_hd__a21o_1 _6142_ (.A1(_2242_),
    .A2(_2960_),
    .B1(_2970_),
    .X(_0425_));
 sky130_fd_sc_hd__buf_6 _6143_ (.A(_2681_),
    .X(_2971_));
 sky130_fd_sc_hd__and3_1 _6144_ (.A(_2971_),
    .B(\dmmu0.page_table[1][8] ),
    .C(_2962_),
    .X(_2972_));
 sky130_fd_sc_hd__a21o_1 _6145_ (.A1(_1946_),
    .A2(_2960_),
    .B1(_2972_),
    .X(_0426_));
 sky130_fd_sc_hd__and3_1 _6146_ (.A(_2971_),
    .B(\dmmu0.page_table[1][9] ),
    .C(_2962_),
    .X(_2973_));
 sky130_fd_sc_hd__a21o_1 _6147_ (.A1(_1948_),
    .A2(_2960_),
    .B1(_2973_),
    .X(_0427_));
 sky130_fd_sc_hd__and3_1 _6148_ (.A(_2971_),
    .B(\dmmu0.page_table[1][10] ),
    .C(_2961_),
    .X(_2974_));
 sky130_fd_sc_hd__a21o_1 _6149_ (.A1(_1950_),
    .A2(_2959_),
    .B1(_2974_),
    .X(_0428_));
 sky130_fd_sc_hd__and3_1 _6150_ (.A(_2971_),
    .B(\dmmu0.page_table[1][11] ),
    .C(_2961_),
    .X(_2975_));
 sky130_fd_sc_hd__a21o_1 _6151_ (.A1(net94),
    .A2(_2959_),
    .B1(_2975_),
    .X(_0429_));
 sky130_fd_sc_hd__and3_1 _6152_ (.A(_2971_),
    .B(\dmmu0.page_table[1][12] ),
    .C(_2961_),
    .X(_2976_));
 sky130_fd_sc_hd__a21o_1 _6153_ (.A1(net95),
    .A2(_2959_),
    .B1(_2976_),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_4 _6154_ (.A(_2931_),
    .X(_2977_));
 sky130_fd_sc_hd__or3_2 _6155_ (.A(net188),
    .B(net181),
    .C(_2062_),
    .X(_2978_));
 sky130_fd_sc_hd__or2_1 _6156_ (.A(_2919_),
    .B(_2978_),
    .X(_2979_));
 sky130_fd_sc_hd__clkbuf_2 _6157_ (.A(_2979_),
    .X(_2980_));
 sky130_fd_sc_hd__clkbuf_4 _6158_ (.A(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__nor2_1 _6159_ (.A(_1968_),
    .B(_2978_),
    .Y(_2982_));
 sky130_fd_sc_hd__buf_2 _6160_ (.A(_2982_),
    .X(_2983_));
 sky130_fd_sc_hd__and2_1 _6161_ (.A(_2879_),
    .B(_2983_),
    .X(_2984_));
 sky130_fd_sc_hd__a31o_1 _6162_ (.A1(_2977_),
    .A2(\dmmu1.page_table[8][0] ),
    .A3(_2981_),
    .B1(_2984_),
    .X(_0431_));
 sky130_fd_sc_hd__and2_1 _6163_ (.A(_2791_),
    .B(_2983_),
    .X(_2985_));
 sky130_fd_sc_hd__a31o_1 _6164_ (.A1(_2977_),
    .A2(\dmmu1.page_table[8][1] ),
    .A3(_2981_),
    .B1(_2985_),
    .X(_0432_));
 sky130_fd_sc_hd__and2_1 _6165_ (.A(_2793_),
    .B(_2983_),
    .X(_2986_));
 sky130_fd_sc_hd__a31o_1 _6166_ (.A1(_2977_),
    .A2(\dmmu1.page_table[8][2] ),
    .A3(_2981_),
    .B1(_2986_),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _6167_ (.A(_2795_),
    .B(_2983_),
    .X(_2987_));
 sky130_fd_sc_hd__a31o_1 _6168_ (.A1(_2977_),
    .A2(\dmmu1.page_table[8][3] ),
    .A3(_2981_),
    .B1(_2987_),
    .X(_0434_));
 sky130_fd_sc_hd__and2_1 _6169_ (.A(_2797_),
    .B(_2983_),
    .X(_2988_));
 sky130_fd_sc_hd__a31o_1 _6170_ (.A1(_2977_),
    .A2(\dmmu1.page_table[8][4] ),
    .A3(_2981_),
    .B1(_2988_),
    .X(_0435_));
 sky130_fd_sc_hd__and2_1 _6171_ (.A(_2799_),
    .B(_2983_),
    .X(_2989_));
 sky130_fd_sc_hd__a31o_1 _6172_ (.A1(_2977_),
    .A2(\dmmu1.page_table[8][5] ),
    .A3(_2981_),
    .B1(_2989_),
    .X(_0436_));
 sky130_fd_sc_hd__and2_1 _6173_ (.A(_2801_),
    .B(_2983_),
    .X(_2990_));
 sky130_fd_sc_hd__a31o_1 _6174_ (.A1(_2977_),
    .A2(\dmmu1.page_table[8][6] ),
    .A3(_2981_),
    .B1(_2990_),
    .X(_0437_));
 sky130_fd_sc_hd__and2_1 _6175_ (.A(_2803_),
    .B(_2983_),
    .X(_2991_));
 sky130_fd_sc_hd__a31o_1 _6176_ (.A1(_2977_),
    .A2(\dmmu1.page_table[8][7] ),
    .A3(_2981_),
    .B1(_2991_),
    .X(_0438_));
 sky130_fd_sc_hd__and2_1 _6177_ (.A(_2891_),
    .B(_2983_),
    .X(_2992_));
 sky130_fd_sc_hd__a31o_1 _6178_ (.A1(_2977_),
    .A2(\dmmu1.page_table[8][8] ),
    .A3(_2981_),
    .B1(_2992_),
    .X(_0439_));
 sky130_fd_sc_hd__and2_1 _6179_ (.A(_2893_),
    .B(_2983_),
    .X(_2993_));
 sky130_fd_sc_hd__a31o_1 _6180_ (.A1(_2977_),
    .A2(\dmmu1.page_table[8][9] ),
    .A3(_2981_),
    .B1(_2993_),
    .X(_0440_));
 sky130_fd_sc_hd__buf_4 _6181_ (.A(_2931_),
    .X(_2994_));
 sky130_fd_sc_hd__and2_1 _6182_ (.A(_2895_),
    .B(_2982_),
    .X(_2995_));
 sky130_fd_sc_hd__a31o_1 _6183_ (.A1(_2994_),
    .A2(\dmmu1.page_table[8][10] ),
    .A3(_2980_),
    .B1(_2995_),
    .X(_0441_));
 sky130_fd_sc_hd__and2_1 _6184_ (.A(_1991_),
    .B(_2982_),
    .X(_2996_));
 sky130_fd_sc_hd__a31o_1 _6185_ (.A1(_2994_),
    .A2(\dmmu1.page_table[8][11] ),
    .A3(_2980_),
    .B1(_2996_),
    .X(_0442_));
 sky130_fd_sc_hd__and2_1 _6186_ (.A(_1993_),
    .B(_2982_),
    .X(_2997_));
 sky130_fd_sc_hd__a31o_1 _6187_ (.A1(_2994_),
    .A2(\dmmu1.page_table[8][12] ),
    .A3(_2980_),
    .B1(_2997_),
    .X(_0443_));
 sky130_fd_sc_hd__or2_1 _6188_ (.A(_2919_),
    .B(_2255_),
    .X(_2998_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _6189_ (.A(_2998_),
    .X(_2999_));
 sky130_fd_sc_hd__buf_4 _6190_ (.A(_2999_),
    .X(_3000_));
 sky130_fd_sc_hd__nor2_1 _6191_ (.A(_1968_),
    .B(_2255_),
    .Y(_3001_));
 sky130_fd_sc_hd__clkbuf_4 _6192_ (.A(_3001_),
    .X(_3002_));
 sky130_fd_sc_hd__and2_1 _6193_ (.A(_2879_),
    .B(_3002_),
    .X(_3003_));
 sky130_fd_sc_hd__a31o_1 _6194_ (.A1(_2994_),
    .A2(\dmmu1.page_table[7][0] ),
    .A3(_3000_),
    .B1(_3003_),
    .X(_0444_));
 sky130_fd_sc_hd__and2_1 _6195_ (.A(_2791_),
    .B(_3002_),
    .X(_3004_));
 sky130_fd_sc_hd__a31o_1 _6196_ (.A1(_2994_),
    .A2(\dmmu1.page_table[7][1] ),
    .A3(_3000_),
    .B1(_3004_),
    .X(_0445_));
 sky130_fd_sc_hd__and2_1 _6197_ (.A(_2793_),
    .B(_3002_),
    .X(_3005_));
 sky130_fd_sc_hd__a31o_1 _6198_ (.A1(_2994_),
    .A2(\dmmu1.page_table[7][2] ),
    .A3(_3000_),
    .B1(_3005_),
    .X(_0446_));
 sky130_fd_sc_hd__and2_1 _6199_ (.A(_2795_),
    .B(_3002_),
    .X(_3006_));
 sky130_fd_sc_hd__a31o_1 _6200_ (.A1(_2994_),
    .A2(\dmmu1.page_table[7][3] ),
    .A3(_3000_),
    .B1(_3006_),
    .X(_0447_));
 sky130_fd_sc_hd__and2_1 _6201_ (.A(_2797_),
    .B(_3002_),
    .X(_3007_));
 sky130_fd_sc_hd__a31o_1 _6202_ (.A1(_2994_),
    .A2(\dmmu1.page_table[7][4] ),
    .A3(_3000_),
    .B1(_3007_),
    .X(_0448_));
 sky130_fd_sc_hd__and2_1 _6203_ (.A(_2799_),
    .B(_3002_),
    .X(_3008_));
 sky130_fd_sc_hd__a31o_1 _6204_ (.A1(_2994_),
    .A2(\dmmu1.page_table[7][5] ),
    .A3(_3000_),
    .B1(_3008_),
    .X(_0449_));
 sky130_fd_sc_hd__and2_1 _6205_ (.A(_2801_),
    .B(_3002_),
    .X(_3009_));
 sky130_fd_sc_hd__a31o_1 _6206_ (.A1(_2994_),
    .A2(\dmmu1.page_table[7][6] ),
    .A3(_3000_),
    .B1(_3009_),
    .X(_0450_));
 sky130_fd_sc_hd__buf_4 _6207_ (.A(_2931_),
    .X(_3010_));
 sky130_fd_sc_hd__and2_1 _6208_ (.A(_2803_),
    .B(_3002_),
    .X(_3011_));
 sky130_fd_sc_hd__a31o_1 _6209_ (.A1(_3010_),
    .A2(\dmmu1.page_table[7][7] ),
    .A3(_3000_),
    .B1(_3011_),
    .X(_0451_));
 sky130_fd_sc_hd__and2_1 _6210_ (.A(_2891_),
    .B(_3002_),
    .X(_3012_));
 sky130_fd_sc_hd__a31o_1 _6211_ (.A1(_3010_),
    .A2(\dmmu1.page_table[7][8] ),
    .A3(_3000_),
    .B1(_3012_),
    .X(_0452_));
 sky130_fd_sc_hd__and2_1 _6212_ (.A(_2893_),
    .B(_3002_),
    .X(_3013_));
 sky130_fd_sc_hd__a31o_1 _6213_ (.A1(_3010_),
    .A2(\dmmu1.page_table[7][9] ),
    .A3(_3000_),
    .B1(_3013_),
    .X(_0453_));
 sky130_fd_sc_hd__and2_1 _6214_ (.A(_2895_),
    .B(_3001_),
    .X(_3014_));
 sky130_fd_sc_hd__a31o_1 _6215_ (.A1(_3010_),
    .A2(\dmmu1.page_table[7][10] ),
    .A3(_2999_),
    .B1(_3014_),
    .X(_0454_));
 sky130_fd_sc_hd__and2_1 _6216_ (.A(_1991_),
    .B(_3001_),
    .X(_3015_));
 sky130_fd_sc_hd__a31o_1 _6217_ (.A1(_3010_),
    .A2(\dmmu1.page_table[7][11] ),
    .A3(_2999_),
    .B1(_3015_),
    .X(_0455_));
 sky130_fd_sc_hd__and2_1 _6218_ (.A(_1993_),
    .B(_3001_),
    .X(_3016_));
 sky130_fd_sc_hd__a31o_1 _6219_ (.A1(_3010_),
    .A2(\dmmu1.page_table[7][12] ),
    .A3(_2999_),
    .B1(_3016_),
    .X(_0456_));
 sky130_fd_sc_hd__or2_1 _6220_ (.A(_2919_),
    .B(_2118_),
    .X(_3017_));
 sky130_fd_sc_hd__clkbuf_2 _6221_ (.A(_3017_),
    .X(_3018_));
 sky130_fd_sc_hd__buf_4 _6222_ (.A(_3018_),
    .X(_3019_));
 sky130_fd_sc_hd__nor2_2 _6223_ (.A(_1968_),
    .B(_2118_),
    .Y(_3020_));
 sky130_fd_sc_hd__clkbuf_4 _6224_ (.A(_3020_),
    .X(_3021_));
 sky130_fd_sc_hd__and2_1 _6225_ (.A(_2879_),
    .B(_3021_),
    .X(_3022_));
 sky130_fd_sc_hd__a31o_1 _6226_ (.A1(_3010_),
    .A2(\dmmu1.page_table[6][0] ),
    .A3(_3019_),
    .B1(_3022_),
    .X(_0457_));
 sky130_fd_sc_hd__and2_1 _6227_ (.A(_2791_),
    .B(_3021_),
    .X(_3023_));
 sky130_fd_sc_hd__a31o_1 _6228_ (.A1(_3010_),
    .A2(\dmmu1.page_table[6][1] ),
    .A3(_3019_),
    .B1(_3023_),
    .X(_0458_));
 sky130_fd_sc_hd__and2_1 _6229_ (.A(_2793_),
    .B(_3021_),
    .X(_3024_));
 sky130_fd_sc_hd__a31o_1 _6230_ (.A1(_3010_),
    .A2(\dmmu1.page_table[6][2] ),
    .A3(_3019_),
    .B1(_3024_),
    .X(_0459_));
 sky130_fd_sc_hd__and2_1 _6231_ (.A(_2795_),
    .B(_3021_),
    .X(_3025_));
 sky130_fd_sc_hd__a31o_1 _6232_ (.A1(_3010_),
    .A2(\dmmu1.page_table[6][3] ),
    .A3(_3019_),
    .B1(_3025_),
    .X(_0460_));
 sky130_fd_sc_hd__buf_4 _6233_ (.A(_2931_),
    .X(_3026_));
 sky130_fd_sc_hd__and2_1 _6234_ (.A(_2797_),
    .B(_3021_),
    .X(_3027_));
 sky130_fd_sc_hd__a31o_1 _6235_ (.A1(_3026_),
    .A2(\dmmu1.page_table[6][4] ),
    .A3(_3019_),
    .B1(_3027_),
    .X(_0461_));
 sky130_fd_sc_hd__and2_1 _6236_ (.A(_2799_),
    .B(_3021_),
    .X(_3028_));
 sky130_fd_sc_hd__a31o_1 _6237_ (.A1(_3026_),
    .A2(\dmmu1.page_table[6][5] ),
    .A3(_3019_),
    .B1(_3028_),
    .X(_0462_));
 sky130_fd_sc_hd__and2_1 _6238_ (.A(_2801_),
    .B(_3021_),
    .X(_3029_));
 sky130_fd_sc_hd__a31o_1 _6239_ (.A1(_3026_),
    .A2(\dmmu1.page_table[6][6] ),
    .A3(_3019_),
    .B1(_3029_),
    .X(_0463_));
 sky130_fd_sc_hd__and2_1 _6240_ (.A(_2803_),
    .B(_3021_),
    .X(_3030_));
 sky130_fd_sc_hd__a31o_1 _6241_ (.A1(_3026_),
    .A2(\dmmu1.page_table[6][7] ),
    .A3(_3019_),
    .B1(_3030_),
    .X(_0464_));
 sky130_fd_sc_hd__and2_1 _6242_ (.A(_2891_),
    .B(_3021_),
    .X(_3031_));
 sky130_fd_sc_hd__a31o_1 _6243_ (.A1(_3026_),
    .A2(\dmmu1.page_table[6][8] ),
    .A3(_3019_),
    .B1(_3031_),
    .X(_0465_));
 sky130_fd_sc_hd__and2_1 _6244_ (.A(_2893_),
    .B(_3021_),
    .X(_3032_));
 sky130_fd_sc_hd__a31o_1 _6245_ (.A1(_3026_),
    .A2(\dmmu1.page_table[6][9] ),
    .A3(_3019_),
    .B1(_3032_),
    .X(_0466_));
 sky130_fd_sc_hd__and2_1 _6246_ (.A(_2895_),
    .B(_3020_),
    .X(_3033_));
 sky130_fd_sc_hd__a31o_1 _6247_ (.A1(_3026_),
    .A2(\dmmu1.page_table[6][10] ),
    .A3(_3018_),
    .B1(_3033_),
    .X(_0467_));
 sky130_fd_sc_hd__and2_1 _6248_ (.A(_1991_),
    .B(_3020_),
    .X(_3034_));
 sky130_fd_sc_hd__a31o_1 _6249_ (.A1(_3026_),
    .A2(\dmmu1.page_table[6][11] ),
    .A3(_3018_),
    .B1(_3034_),
    .X(_0468_));
 sky130_fd_sc_hd__and2_1 _6250_ (.A(_1993_),
    .B(_3020_),
    .X(_3035_));
 sky130_fd_sc_hd__a31o_1 _6251_ (.A1(_3026_),
    .A2(\dmmu1.page_table[6][12] ),
    .A3(_3018_),
    .B1(_3035_),
    .X(_0469_));
 sky130_fd_sc_hd__or2_1 _6252_ (.A(_2919_),
    .B(_2136_),
    .X(_3036_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _6253_ (.A(_3036_),
    .X(_3037_));
 sky130_fd_sc_hd__buf_4 _6254_ (.A(_3037_),
    .X(_3038_));
 sky130_fd_sc_hd__nor2_1 _6255_ (.A(_2784_),
    .B(_2136_),
    .Y(_3039_));
 sky130_fd_sc_hd__clkbuf_4 _6256_ (.A(_3039_),
    .X(_3040_));
 sky130_fd_sc_hd__and2_1 _6257_ (.A(_2879_),
    .B(_3040_),
    .X(_3041_));
 sky130_fd_sc_hd__a31o_1 _6258_ (.A1(_3026_),
    .A2(\dmmu1.page_table[5][0] ),
    .A3(_3038_),
    .B1(_3041_),
    .X(_0470_));
 sky130_fd_sc_hd__buf_4 _6259_ (.A(_2931_),
    .X(_3042_));
 sky130_fd_sc_hd__and2_1 _6260_ (.A(_2791_),
    .B(_3040_),
    .X(_3043_));
 sky130_fd_sc_hd__a31o_1 _6261_ (.A1(_3042_),
    .A2(\dmmu1.page_table[5][1] ),
    .A3(_3038_),
    .B1(_3043_),
    .X(_0471_));
 sky130_fd_sc_hd__and2_1 _6262_ (.A(_2793_),
    .B(_3040_),
    .X(_3044_));
 sky130_fd_sc_hd__a31o_1 _6263_ (.A1(_3042_),
    .A2(\dmmu1.page_table[5][2] ),
    .A3(_3038_),
    .B1(_3044_),
    .X(_0472_));
 sky130_fd_sc_hd__and2_1 _6264_ (.A(_2795_),
    .B(_3040_),
    .X(_3045_));
 sky130_fd_sc_hd__a31o_1 _6265_ (.A1(_3042_),
    .A2(\dmmu1.page_table[5][3] ),
    .A3(_3038_),
    .B1(_3045_),
    .X(_0473_));
 sky130_fd_sc_hd__and2_1 _6266_ (.A(_2797_),
    .B(_3040_),
    .X(_3046_));
 sky130_fd_sc_hd__a31o_1 _6267_ (.A1(_3042_),
    .A2(\dmmu1.page_table[5][4] ),
    .A3(_3038_),
    .B1(_3046_),
    .X(_0474_));
 sky130_fd_sc_hd__and2_1 _6268_ (.A(_2799_),
    .B(_3040_),
    .X(_3047_));
 sky130_fd_sc_hd__a31o_1 _6269_ (.A1(_3042_),
    .A2(\dmmu1.page_table[5][5] ),
    .A3(_3038_),
    .B1(_3047_),
    .X(_0475_));
 sky130_fd_sc_hd__and2_1 _6270_ (.A(_2801_),
    .B(_3040_),
    .X(_3048_));
 sky130_fd_sc_hd__a31o_1 _6271_ (.A1(_3042_),
    .A2(\dmmu1.page_table[5][6] ),
    .A3(_3038_),
    .B1(_3048_),
    .X(_0476_));
 sky130_fd_sc_hd__and2_1 _6272_ (.A(_2803_),
    .B(_3040_),
    .X(_3049_));
 sky130_fd_sc_hd__a31o_1 _6273_ (.A1(_3042_),
    .A2(\dmmu1.page_table[5][7] ),
    .A3(_3038_),
    .B1(_3049_),
    .X(_0477_));
 sky130_fd_sc_hd__and2_1 _6274_ (.A(_2891_),
    .B(_3040_),
    .X(_3050_));
 sky130_fd_sc_hd__a31o_1 _6275_ (.A1(_3042_),
    .A2(\dmmu1.page_table[5][8] ),
    .A3(_3038_),
    .B1(_3050_),
    .X(_0478_));
 sky130_fd_sc_hd__and2_1 _6276_ (.A(_2893_),
    .B(_3040_),
    .X(_3051_));
 sky130_fd_sc_hd__a31o_1 _6277_ (.A1(_3042_),
    .A2(\dmmu1.page_table[5][9] ),
    .A3(_3038_),
    .B1(_3051_),
    .X(_0479_));
 sky130_fd_sc_hd__and2_1 _6278_ (.A(_2895_),
    .B(_3039_),
    .X(_3052_));
 sky130_fd_sc_hd__a31o_1 _6279_ (.A1(_3042_),
    .A2(\dmmu1.page_table[5][10] ),
    .A3(_3037_),
    .B1(_3052_),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_4 _6280_ (.A(_2931_),
    .X(_3053_));
 sky130_fd_sc_hd__and2_1 _6281_ (.A(net199),
    .B(_3039_),
    .X(_3054_));
 sky130_fd_sc_hd__a31o_1 _6282_ (.A1(_3053_),
    .A2(\dmmu1.page_table[5][11] ),
    .A3(_3037_),
    .B1(_3054_),
    .X(_0481_));
 sky130_fd_sc_hd__and2_1 _6283_ (.A(net200),
    .B(_3039_),
    .X(_3055_));
 sky130_fd_sc_hd__a31o_1 _6284_ (.A1(_3053_),
    .A2(\dmmu1.page_table[5][12] ),
    .A3(_3037_),
    .B1(_3055_),
    .X(_0482_));
 sky130_fd_sc_hd__or2_1 _6285_ (.A(_2919_),
    .B(_2153_),
    .X(_3056_));
 sky130_fd_sc_hd__clkbuf_2 _6286_ (.A(_3056_),
    .X(_3057_));
 sky130_fd_sc_hd__clkbuf_4 _6287_ (.A(_3057_),
    .X(_3058_));
 sky130_fd_sc_hd__nor2_2 _6288_ (.A(_2784_),
    .B(_2153_),
    .Y(_3059_));
 sky130_fd_sc_hd__buf_2 _6289_ (.A(_3059_),
    .X(_3060_));
 sky130_fd_sc_hd__and2_1 _6290_ (.A(_2879_),
    .B(_3060_),
    .X(_3061_));
 sky130_fd_sc_hd__a31o_1 _6291_ (.A1(_3053_),
    .A2(\dmmu1.page_table[4][0] ),
    .A3(_3058_),
    .B1(_3061_),
    .X(_0483_));
 sky130_fd_sc_hd__and2_1 _6292_ (.A(net201),
    .B(_3060_),
    .X(_3062_));
 sky130_fd_sc_hd__a31o_1 _6293_ (.A1(_3053_),
    .A2(\dmmu1.page_table[4][1] ),
    .A3(_3058_),
    .B1(_3062_),
    .X(_0484_));
 sky130_fd_sc_hd__and2_1 _6294_ (.A(net202),
    .B(_3060_),
    .X(_3063_));
 sky130_fd_sc_hd__a31o_1 _6295_ (.A1(_3053_),
    .A2(\dmmu1.page_table[4][2] ),
    .A3(_3058_),
    .B1(_3063_),
    .X(_0485_));
 sky130_fd_sc_hd__and2_1 _6296_ (.A(net203),
    .B(_3060_),
    .X(_3064_));
 sky130_fd_sc_hd__a31o_1 _6297_ (.A1(_3053_),
    .A2(\dmmu1.page_table[4][3] ),
    .A3(_3058_),
    .B1(_3064_),
    .X(_0486_));
 sky130_fd_sc_hd__and2_1 _6298_ (.A(net204),
    .B(_3060_),
    .X(_3065_));
 sky130_fd_sc_hd__a31o_1 _6299_ (.A1(_3053_),
    .A2(\dmmu1.page_table[4][4] ),
    .A3(_3058_),
    .B1(_3065_),
    .X(_0487_));
 sky130_fd_sc_hd__and2_1 _6300_ (.A(net205),
    .B(_3060_),
    .X(_3066_));
 sky130_fd_sc_hd__a31o_1 _6301_ (.A1(_3053_),
    .A2(\dmmu1.page_table[4][5] ),
    .A3(_3058_),
    .B1(_3066_),
    .X(_0488_));
 sky130_fd_sc_hd__and2_1 _6302_ (.A(net206),
    .B(_3060_),
    .X(_3067_));
 sky130_fd_sc_hd__a31o_1 _6303_ (.A1(_3053_),
    .A2(\dmmu1.page_table[4][6] ),
    .A3(_3058_),
    .B1(_3067_),
    .X(_0489_));
 sky130_fd_sc_hd__and2_1 _6304_ (.A(net207),
    .B(_3060_),
    .X(_3068_));
 sky130_fd_sc_hd__a31o_1 _6305_ (.A1(_3053_),
    .A2(\dmmu1.page_table[4][7] ),
    .A3(_3058_),
    .B1(_3068_),
    .X(_0490_));
 sky130_fd_sc_hd__buf_4 _6306_ (.A(_2931_),
    .X(_3069_));
 sky130_fd_sc_hd__and2_1 _6307_ (.A(_2891_),
    .B(_3060_),
    .X(_3070_));
 sky130_fd_sc_hd__a31o_1 _6308_ (.A1(_3069_),
    .A2(\dmmu1.page_table[4][8] ),
    .A3(_3058_),
    .B1(_3070_),
    .X(_0491_));
 sky130_fd_sc_hd__and2_1 _6309_ (.A(_2893_),
    .B(_3060_),
    .X(_3071_));
 sky130_fd_sc_hd__a31o_1 _6310_ (.A1(_3069_),
    .A2(\dmmu1.page_table[4][9] ),
    .A3(_3058_),
    .B1(_3071_),
    .X(_0492_));
 sky130_fd_sc_hd__and2_1 _6311_ (.A(_2895_),
    .B(_3059_),
    .X(_3072_));
 sky130_fd_sc_hd__a31o_1 _6312_ (.A1(_3069_),
    .A2(\dmmu1.page_table[4][10] ),
    .A3(_3057_),
    .B1(_3072_),
    .X(_0493_));
 sky130_fd_sc_hd__and2_1 _6313_ (.A(net199),
    .B(_3059_),
    .X(_3073_));
 sky130_fd_sc_hd__a31o_1 _6314_ (.A1(_3069_),
    .A2(\dmmu1.page_table[4][11] ),
    .A3(_3057_),
    .B1(_3073_),
    .X(_0494_));
 sky130_fd_sc_hd__and2_1 _6315_ (.A(net200),
    .B(_3059_),
    .X(_3074_));
 sky130_fd_sc_hd__a31o_1 _6316_ (.A1(_3069_),
    .A2(\dmmu1.page_table[4][12] ),
    .A3(_3057_),
    .B1(_3074_),
    .X(_0495_));
 sky130_fd_sc_hd__or2_1 _6317_ (.A(_2919_),
    .B(_2193_),
    .X(_3075_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _6318_ (.A(_3075_),
    .X(_3076_));
 sky130_fd_sc_hd__clkbuf_4 _6319_ (.A(_3076_),
    .X(_3077_));
 sky130_fd_sc_hd__nor2_1 _6320_ (.A(_2784_),
    .B(_2193_),
    .Y(_3078_));
 sky130_fd_sc_hd__clkbuf_4 _6321_ (.A(_3078_),
    .X(_3079_));
 sky130_fd_sc_hd__and2_1 _6322_ (.A(_2879_),
    .B(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__a31o_1 _6323_ (.A1(_3069_),
    .A2(\dmmu1.page_table[3][0] ),
    .A3(_3077_),
    .B1(_3080_),
    .X(_0496_));
 sky130_fd_sc_hd__and2_1 _6324_ (.A(net201),
    .B(_3079_),
    .X(_3081_));
 sky130_fd_sc_hd__a31o_1 _6325_ (.A1(_3069_),
    .A2(\dmmu1.page_table[3][1] ),
    .A3(_3077_),
    .B1(_3081_),
    .X(_0497_));
 sky130_fd_sc_hd__and2_1 _6326_ (.A(net202),
    .B(_3079_),
    .X(_3082_));
 sky130_fd_sc_hd__a31o_1 _6327_ (.A1(_3069_),
    .A2(\dmmu1.page_table[3][2] ),
    .A3(_3077_),
    .B1(_3082_),
    .X(_0498_));
 sky130_fd_sc_hd__and2_1 _6328_ (.A(net203),
    .B(_3079_),
    .X(_3083_));
 sky130_fd_sc_hd__a31o_1 _6329_ (.A1(_3069_),
    .A2(\dmmu1.page_table[3][3] ),
    .A3(_3077_),
    .B1(_3083_),
    .X(_0499_));
 sky130_fd_sc_hd__and2_1 _6330_ (.A(net204),
    .B(_3079_),
    .X(_3084_));
 sky130_fd_sc_hd__a31o_1 _6331_ (.A1(_3069_),
    .A2(\dmmu1.page_table[3][4] ),
    .A3(_3077_),
    .B1(_3084_),
    .X(_0500_));
 sky130_fd_sc_hd__buf_4 _6332_ (.A(_2931_),
    .X(_3085_));
 sky130_fd_sc_hd__and2_1 _6333_ (.A(net205),
    .B(_3079_),
    .X(_3086_));
 sky130_fd_sc_hd__a31o_1 _6334_ (.A1(_3085_),
    .A2(\dmmu1.page_table[3][5] ),
    .A3(_3077_),
    .B1(_3086_),
    .X(_0501_));
 sky130_fd_sc_hd__and2_1 _6335_ (.A(net206),
    .B(_3079_),
    .X(_3087_));
 sky130_fd_sc_hd__a31o_1 _6336_ (.A1(_3085_),
    .A2(\dmmu1.page_table[3][6] ),
    .A3(_3077_),
    .B1(_3087_),
    .X(_0502_));
 sky130_fd_sc_hd__and2_1 _6337_ (.A(net207),
    .B(_3079_),
    .X(_3088_));
 sky130_fd_sc_hd__a31o_1 _6338_ (.A1(_3085_),
    .A2(\dmmu1.page_table[3][7] ),
    .A3(_3077_),
    .B1(_3088_),
    .X(_0503_));
 sky130_fd_sc_hd__and2_1 _6339_ (.A(_2891_),
    .B(_3079_),
    .X(_3089_));
 sky130_fd_sc_hd__a31o_1 _6340_ (.A1(_3085_),
    .A2(\dmmu1.page_table[3][8] ),
    .A3(_3077_),
    .B1(_3089_),
    .X(_0504_));
 sky130_fd_sc_hd__and2_1 _6341_ (.A(_2893_),
    .B(_3079_),
    .X(_3090_));
 sky130_fd_sc_hd__a31o_1 _6342_ (.A1(_3085_),
    .A2(\dmmu1.page_table[3][9] ),
    .A3(_3077_),
    .B1(_3090_),
    .X(_0505_));
 sky130_fd_sc_hd__and2_1 _6343_ (.A(_2895_),
    .B(_3078_),
    .X(_3091_));
 sky130_fd_sc_hd__a31o_1 _6344_ (.A1(_3085_),
    .A2(\dmmu1.page_table[3][10] ),
    .A3(_3076_),
    .B1(_3091_),
    .X(_0506_));
 sky130_fd_sc_hd__and2_1 _6345_ (.A(net199),
    .B(_3078_),
    .X(_3092_));
 sky130_fd_sc_hd__a31o_1 _6346_ (.A1(_3085_),
    .A2(\dmmu1.page_table[3][11] ),
    .A3(_3076_),
    .B1(_3092_),
    .X(_0507_));
 sky130_fd_sc_hd__and2_1 _6347_ (.A(net200),
    .B(_3078_),
    .X(_3093_));
 sky130_fd_sc_hd__a31o_1 _6348_ (.A1(_3085_),
    .A2(\dmmu1.page_table[3][12] ),
    .A3(_3076_),
    .B1(_3093_),
    .X(_0508_));
 sky130_fd_sc_hd__or2_1 _6349_ (.A(_2919_),
    .B(_2170_),
    .X(_3094_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _6350_ (.A(_3094_),
    .X(_3095_));
 sky130_fd_sc_hd__clkbuf_4 _6351_ (.A(_3095_),
    .X(_3096_));
 sky130_fd_sc_hd__nor2_1 _6352_ (.A(_2784_),
    .B(_2170_),
    .Y(_3097_));
 sky130_fd_sc_hd__buf_2 _6353_ (.A(_3097_),
    .X(_3098_));
 sky130_fd_sc_hd__and2_1 _6354_ (.A(net197),
    .B(_3098_),
    .X(_3099_));
 sky130_fd_sc_hd__a31o_1 _6355_ (.A1(_3085_),
    .A2(\dmmu1.page_table[2][0] ),
    .A3(_3096_),
    .B1(_3099_),
    .X(_0509_));
 sky130_fd_sc_hd__and2_1 _6356_ (.A(net201),
    .B(_3098_),
    .X(_3100_));
 sky130_fd_sc_hd__a31o_1 _6357_ (.A1(_3085_),
    .A2(\dmmu1.page_table[2][1] ),
    .A3(_3096_),
    .B1(_3100_),
    .X(_0510_));
 sky130_fd_sc_hd__clkbuf_4 _6358_ (.A(_1910_),
    .X(_3101_));
 sky130_fd_sc_hd__and2_1 _6359_ (.A(net202),
    .B(_3098_),
    .X(_3102_));
 sky130_fd_sc_hd__a31o_1 _6360_ (.A1(_3101_),
    .A2(\dmmu1.page_table[2][2] ),
    .A3(_3096_),
    .B1(_3102_),
    .X(_0511_));
 sky130_fd_sc_hd__and2_1 _6361_ (.A(net203),
    .B(_3098_),
    .X(_3103_));
 sky130_fd_sc_hd__a31o_1 _6362_ (.A1(_3101_),
    .A2(\dmmu1.page_table[2][3] ),
    .A3(_3096_),
    .B1(_3103_),
    .X(_0512_));
 sky130_fd_sc_hd__and2_1 _6363_ (.A(net204),
    .B(_3098_),
    .X(_3104_));
 sky130_fd_sc_hd__a31o_1 _6364_ (.A1(_3101_),
    .A2(\dmmu1.page_table[2][4] ),
    .A3(_3096_),
    .B1(_3104_),
    .X(_0513_));
 sky130_fd_sc_hd__and2_1 _6365_ (.A(net205),
    .B(_3098_),
    .X(_3105_));
 sky130_fd_sc_hd__a31o_1 _6366_ (.A1(_3101_),
    .A2(\dmmu1.page_table[2][5] ),
    .A3(_3096_),
    .B1(_3105_),
    .X(_0514_));
 sky130_fd_sc_hd__and2_1 _6367_ (.A(net206),
    .B(_3098_),
    .X(_3106_));
 sky130_fd_sc_hd__a31o_1 _6368_ (.A1(_3101_),
    .A2(\dmmu1.page_table[2][6] ),
    .A3(_3096_),
    .B1(_3106_),
    .X(_0515_));
 sky130_fd_sc_hd__and2_1 _6369_ (.A(net207),
    .B(_3098_),
    .X(_3107_));
 sky130_fd_sc_hd__a31o_1 _6370_ (.A1(_3101_),
    .A2(\dmmu1.page_table[2][7] ),
    .A3(_3096_),
    .B1(_3107_),
    .X(_0516_));
 sky130_fd_sc_hd__and2_1 _6371_ (.A(net208),
    .B(_3098_),
    .X(_3108_));
 sky130_fd_sc_hd__a31o_1 _6372_ (.A1(_3101_),
    .A2(\dmmu1.page_table[2][8] ),
    .A3(_3096_),
    .B1(_3108_),
    .X(_0517_));
 sky130_fd_sc_hd__and2_1 _6373_ (.A(net209),
    .B(_3098_),
    .X(_3109_));
 sky130_fd_sc_hd__a31o_1 _6374_ (.A1(_3101_),
    .A2(\dmmu1.page_table[2][9] ),
    .A3(_3096_),
    .B1(_3109_),
    .X(_0518_));
 sky130_fd_sc_hd__and2_1 _6375_ (.A(net198),
    .B(_3097_),
    .X(_3110_));
 sky130_fd_sc_hd__a31o_1 _6376_ (.A1(_3101_),
    .A2(\dmmu1.page_table[2][10] ),
    .A3(_3095_),
    .B1(_3110_),
    .X(_0519_));
 sky130_fd_sc_hd__and2_1 _6377_ (.A(net199),
    .B(_3097_),
    .X(_3111_));
 sky130_fd_sc_hd__a31o_1 _6378_ (.A1(_3101_),
    .A2(\dmmu1.page_table[2][11] ),
    .A3(_3095_),
    .B1(_3111_),
    .X(_0520_));
 sky130_fd_sc_hd__clkbuf_4 _6379_ (.A(_1910_),
    .X(_3112_));
 sky130_fd_sc_hd__and2_1 _6380_ (.A(net200),
    .B(_3097_),
    .X(_3113_));
 sky130_fd_sc_hd__a31o_1 _6381_ (.A1(_3112_),
    .A2(\dmmu1.page_table[2][12] ),
    .A3(_3095_),
    .B1(_3113_),
    .X(_0521_));
 sky130_fd_sc_hd__or2_1 _6382_ (.A(_2919_),
    .B(_2187_),
    .X(_3114_));
 sky130_fd_sc_hd__clkbuf_2 _6383_ (.A(_3114_),
    .X(_3115_));
 sky130_fd_sc_hd__clkbuf_4 _6384_ (.A(_3115_),
    .X(_3116_));
 sky130_fd_sc_hd__nor2_1 _6385_ (.A(_2784_),
    .B(_2187_),
    .Y(_3117_));
 sky130_fd_sc_hd__buf_2 _6386_ (.A(_3117_),
    .X(_3118_));
 sky130_fd_sc_hd__and2_1 _6387_ (.A(net197),
    .B(_3118_),
    .X(_3119_));
 sky130_fd_sc_hd__a31o_1 _6388_ (.A1(_3112_),
    .A2(\dmmu1.page_table[1][0] ),
    .A3(_3116_),
    .B1(_3119_),
    .X(_0522_));
 sky130_fd_sc_hd__and2_1 _6389_ (.A(net201),
    .B(_3118_),
    .X(_3120_));
 sky130_fd_sc_hd__a31o_1 _6390_ (.A1(_3112_),
    .A2(\dmmu1.page_table[1][1] ),
    .A3(_3116_),
    .B1(_3120_),
    .X(_0523_));
 sky130_fd_sc_hd__and2_1 _6391_ (.A(net202),
    .B(_3118_),
    .X(_3121_));
 sky130_fd_sc_hd__a31o_1 _6392_ (.A1(_3112_),
    .A2(\dmmu1.page_table[1][2] ),
    .A3(_3116_),
    .B1(_3121_),
    .X(_0524_));
 sky130_fd_sc_hd__and2_1 _6393_ (.A(net203),
    .B(_3118_),
    .X(_3122_));
 sky130_fd_sc_hd__a31o_1 _6394_ (.A1(_3112_),
    .A2(\dmmu1.page_table[1][3] ),
    .A3(_3116_),
    .B1(_3122_),
    .X(_0525_));
 sky130_fd_sc_hd__and2_1 _6395_ (.A(net204),
    .B(_3118_),
    .X(_3123_));
 sky130_fd_sc_hd__a31o_1 _6396_ (.A1(_3112_),
    .A2(\dmmu1.page_table[1][4] ),
    .A3(_3116_),
    .B1(_3123_),
    .X(_0526_));
 sky130_fd_sc_hd__and2_1 _6397_ (.A(net205),
    .B(_3118_),
    .X(_3124_));
 sky130_fd_sc_hd__a31o_1 _6398_ (.A1(_3112_),
    .A2(\dmmu1.page_table[1][5] ),
    .A3(_3116_),
    .B1(_3124_),
    .X(_0527_));
 sky130_fd_sc_hd__and2_1 _6399_ (.A(net206),
    .B(_3118_),
    .X(_3125_));
 sky130_fd_sc_hd__a31o_1 _6400_ (.A1(_3112_),
    .A2(\dmmu1.page_table[1][6] ),
    .A3(_3116_),
    .B1(_3125_),
    .X(_0528_));
 sky130_fd_sc_hd__and2_1 _6401_ (.A(net207),
    .B(_3118_),
    .X(_3126_));
 sky130_fd_sc_hd__a31o_1 _6402_ (.A1(_3112_),
    .A2(\dmmu1.page_table[1][7] ),
    .A3(_3116_),
    .B1(_3126_),
    .X(_0529_));
 sky130_fd_sc_hd__and2_1 _6403_ (.A(net208),
    .B(_3118_),
    .X(_3127_));
 sky130_fd_sc_hd__a31o_1 _6404_ (.A1(_3112_),
    .A2(\dmmu1.page_table[1][8] ),
    .A3(_3116_),
    .B1(_3127_),
    .X(_0530_));
 sky130_fd_sc_hd__buf_4 _6405_ (.A(_1910_),
    .X(_3128_));
 sky130_fd_sc_hd__and2_1 _6406_ (.A(net209),
    .B(_3118_),
    .X(_3129_));
 sky130_fd_sc_hd__a31o_1 _6407_ (.A1(_3128_),
    .A2(\dmmu1.page_table[1][9] ),
    .A3(_3116_),
    .B1(_3129_),
    .X(_0531_));
 sky130_fd_sc_hd__and2_1 _6408_ (.A(net198),
    .B(_3117_),
    .X(_3130_));
 sky130_fd_sc_hd__a31o_1 _6409_ (.A1(_3128_),
    .A2(\dmmu1.page_table[1][10] ),
    .A3(_3115_),
    .B1(_3130_),
    .X(_0532_));
 sky130_fd_sc_hd__and2_1 _6410_ (.A(net199),
    .B(_3117_),
    .X(_3131_));
 sky130_fd_sc_hd__a31o_1 _6411_ (.A1(_3128_),
    .A2(\dmmu1.page_table[1][11] ),
    .A3(_3115_),
    .B1(_3131_),
    .X(_0533_));
 sky130_fd_sc_hd__and2_1 _6412_ (.A(net200),
    .B(_3117_),
    .X(_3132_));
 sky130_fd_sc_hd__a31o_1 _6413_ (.A1(_3128_),
    .A2(\dmmu1.page_table[1][12] ),
    .A3(_3115_),
    .B1(_3132_),
    .X(_0534_));
 sky130_fd_sc_hd__or2_1 _6414_ (.A(_1958_),
    .B(_2272_),
    .X(_3133_));
 sky130_fd_sc_hd__clkbuf_2 _6415_ (.A(_3133_),
    .X(_3134_));
 sky130_fd_sc_hd__clkbuf_4 _6416_ (.A(_3134_),
    .X(_3135_));
 sky130_fd_sc_hd__nor2_1 _6417_ (.A(_2784_),
    .B(_2272_),
    .Y(_3136_));
 sky130_fd_sc_hd__buf_2 _6418_ (.A(_3136_),
    .X(_3137_));
 sky130_fd_sc_hd__and2_1 _6419_ (.A(net197),
    .B(_3137_),
    .X(_3138_));
 sky130_fd_sc_hd__a31o_1 _6420_ (.A1(_3128_),
    .A2(\dmmu1.page_table[0][0] ),
    .A3(_3135_),
    .B1(_3138_),
    .X(_0535_));
 sky130_fd_sc_hd__and2_1 _6421_ (.A(net201),
    .B(_3137_),
    .X(_3139_));
 sky130_fd_sc_hd__a31o_1 _6422_ (.A1(_3128_),
    .A2(\dmmu1.page_table[0][1] ),
    .A3(_3135_),
    .B1(_3139_),
    .X(_0536_));
 sky130_fd_sc_hd__and2_1 _6423_ (.A(net202),
    .B(_3137_),
    .X(_3140_));
 sky130_fd_sc_hd__a31o_1 _6424_ (.A1(_3128_),
    .A2(\dmmu1.page_table[0][2] ),
    .A3(_3135_),
    .B1(_3140_),
    .X(_0537_));
 sky130_fd_sc_hd__and2_1 _6425_ (.A(net203),
    .B(_3137_),
    .X(_3141_));
 sky130_fd_sc_hd__a31o_1 _6426_ (.A1(_3128_),
    .A2(\dmmu1.page_table[0][3] ),
    .A3(_3135_),
    .B1(_3141_),
    .X(_0538_));
 sky130_fd_sc_hd__and2_1 _6427_ (.A(net204),
    .B(_3137_),
    .X(_3142_));
 sky130_fd_sc_hd__a31o_1 _6428_ (.A1(_3128_),
    .A2(\dmmu1.page_table[0][4] ),
    .A3(_3135_),
    .B1(_3142_),
    .X(_0539_));
 sky130_fd_sc_hd__and2_1 _6429_ (.A(net205),
    .B(_3137_),
    .X(_3143_));
 sky130_fd_sc_hd__a31o_1 _6430_ (.A1(_3128_),
    .A2(\dmmu1.page_table[0][5] ),
    .A3(_3135_),
    .B1(_3143_),
    .X(_0540_));
 sky130_fd_sc_hd__and2_1 _6431_ (.A(net206),
    .B(_3137_),
    .X(_3144_));
 sky130_fd_sc_hd__a31o_1 _6432_ (.A1(_1898_),
    .A2(\dmmu1.page_table[0][6] ),
    .A3(_3135_),
    .B1(_3144_),
    .X(_0541_));
 sky130_fd_sc_hd__and2_1 _6433_ (.A(net207),
    .B(_3137_),
    .X(_3145_));
 sky130_fd_sc_hd__a31o_1 _6434_ (.A1(_1898_),
    .A2(\dmmu1.page_table[0][7] ),
    .A3(_3135_),
    .B1(_3145_),
    .X(_0542_));
 sky130_fd_sc_hd__and2_1 _6435_ (.A(net208),
    .B(_3137_),
    .X(_3146_));
 sky130_fd_sc_hd__a31o_1 _6436_ (.A1(_1898_),
    .A2(\dmmu1.page_table[0][8] ),
    .A3(_3135_),
    .B1(_3146_),
    .X(_0543_));
 sky130_fd_sc_hd__and2_1 _6437_ (.A(net209),
    .B(_3137_),
    .X(_3147_));
 sky130_fd_sc_hd__a31o_1 _6438_ (.A1(_1898_),
    .A2(\dmmu1.page_table[0][9] ),
    .A3(_3135_),
    .B1(_3147_),
    .X(_0544_));
 sky130_fd_sc_hd__and2_1 _6439_ (.A(net198),
    .B(_3136_),
    .X(_3148_));
 sky130_fd_sc_hd__a31o_1 _6440_ (.A1(_1898_),
    .A2(\dmmu1.page_table[0][10] ),
    .A3(_3134_),
    .B1(_3148_),
    .X(_0545_));
 sky130_fd_sc_hd__and2_1 _6441_ (.A(net199),
    .B(_3136_),
    .X(_3149_));
 sky130_fd_sc_hd__a31o_1 _6442_ (.A1(_1898_),
    .A2(\dmmu1.page_table[0][11] ),
    .A3(_3134_),
    .B1(_3149_),
    .X(_0546_));
 sky130_fd_sc_hd__and2_1 _6443_ (.A(net200),
    .B(_3136_),
    .X(_3150_));
 sky130_fd_sc_hd__a31o_1 _6444_ (.A1(_1898_),
    .A2(\dmmu1.page_table[0][12] ),
    .A3(_3134_),
    .B1(_3150_),
    .X(_0547_));
 sky130_fd_sc_hd__nor2_1 _6445_ (.A(net213),
    .B(net212),
    .Y(_3151_));
 sky130_fd_sc_hd__a21o_1 _6446_ (.A1(net562),
    .A2(_3151_),
    .B1(\mem_dcache_arb.select ),
    .X(_3152_));
 sky130_fd_sc_hd__o311a_1 _6447_ (.A1(net213),
    .A2(net212),
    .A3(_0817_),
    .B1(_3152_),
    .C1(_1911_),
    .X(_0548_));
 sky130_fd_sc_hd__nor3_1 _6448_ (.A(net211),
    .B(_0810_),
    .C(_0819_),
    .Y(_0549_));
 sky130_fd_sc_hd__inv_2 _6449_ (.A(\mem_dcache_arb.transfer_active ),
    .Y(_3153_));
 sky130_fd_sc_hd__nor2_1 _6450_ (.A(net710),
    .B(_0809_),
    .Y(_3154_));
 sky130_fd_sc_hd__o211a_1 _6451_ (.A1(_3153_),
    .A2(\mem_dcache_arb.select ),
    .B1(_0817_),
    .C1(_3154_),
    .X(_0550_));
 sky130_fd_sc_hd__a311o_1 _6452_ (.A1(_3153_),
    .A2(_0809_),
    .A3(_0810_),
    .B1(net213),
    .C1(net212),
    .X(_3155_));
 sky130_fd_sc_hd__nor2_1 _6453_ (.A(net710),
    .B(_3155_),
    .Y(_0551_));
 sky130_fd_sc_hd__nor2_1 _6454_ (.A(_1999_),
    .B(_2978_),
    .Y(_3156_));
 sky130_fd_sc_hd__clkbuf_4 _6455_ (.A(_3156_),
    .X(_3157_));
 sky130_fd_sc_hd__or2_1 _6456_ (.A(_2084_),
    .B(_2978_),
    .X(_3158_));
 sky130_fd_sc_hd__buf_2 _6457_ (.A(_3158_),
    .X(_3159_));
 sky130_fd_sc_hd__and3_1 _6458_ (.A(_2971_),
    .B(\immu_1.page_table[8][0] ),
    .C(_3159_),
    .X(_3160_));
 sky130_fd_sc_hd__a21o_1 _6459_ (.A1(_1995_),
    .A2(_3157_),
    .B1(_3160_),
    .X(_0552_));
 sky130_fd_sc_hd__and3_1 _6460_ (.A(_2971_),
    .B(\immu_1.page_table[8][1] ),
    .C(_3159_),
    .X(_3161_));
 sky130_fd_sc_hd__a21o_1 _6461_ (.A1(_1967_),
    .A2(_3157_),
    .B1(_3161_),
    .X(_0553_));
 sky130_fd_sc_hd__and3_1 _6462_ (.A(_2971_),
    .B(\immu_1.page_table[8][2] ),
    .C(_3159_),
    .X(_3162_));
 sky130_fd_sc_hd__a21o_1 _6463_ (.A1(_1972_),
    .A2(_3157_),
    .B1(_3162_),
    .X(_0554_));
 sky130_fd_sc_hd__and3_1 _6464_ (.A(_2971_),
    .B(\immu_1.page_table[8][3] ),
    .C(_3159_),
    .X(_3163_));
 sky130_fd_sc_hd__a21o_1 _6465_ (.A1(_1974_),
    .A2(_3157_),
    .B1(_3163_),
    .X(_0555_));
 sky130_fd_sc_hd__and3_1 _6466_ (.A(_2971_),
    .B(\immu_1.page_table[8][4] ),
    .C(_3159_),
    .X(_3164_));
 sky130_fd_sc_hd__a21o_1 _6467_ (.A1(_1977_),
    .A2(_3157_),
    .B1(_3164_),
    .X(_0556_));
 sky130_fd_sc_hd__and3_1 _6468_ (.A(_2190_),
    .B(\immu_1.page_table[8][5] ),
    .C(_3159_),
    .X(_3165_));
 sky130_fd_sc_hd__a21o_1 _6469_ (.A1(_1979_),
    .A2(_3157_),
    .B1(_3165_),
    .X(_0557_));
 sky130_fd_sc_hd__and3_1 _6470_ (.A(_2190_),
    .B(\immu_1.page_table[8][6] ),
    .C(_3159_),
    .X(_3166_));
 sky130_fd_sc_hd__a21o_1 _6471_ (.A1(_1981_),
    .A2(_3157_),
    .B1(_3166_),
    .X(_0558_));
 sky130_fd_sc_hd__and3_1 _6472_ (.A(_2190_),
    .B(\immu_1.page_table[8][7] ),
    .C(_3159_),
    .X(_3167_));
 sky130_fd_sc_hd__a21o_1 _6473_ (.A1(_1983_),
    .A2(_3157_),
    .B1(_3167_),
    .X(_0559_));
 sky130_fd_sc_hd__and3_1 _6474_ (.A(_2190_),
    .B(\immu_1.page_table[8][8] ),
    .C(_3159_),
    .X(_3168_));
 sky130_fd_sc_hd__a21o_1 _6475_ (.A1(_1985_),
    .A2(_3157_),
    .B1(_3168_),
    .X(_0560_));
 sky130_fd_sc_hd__and3_1 _6476_ (.A(_2190_),
    .B(\immu_1.page_table[8][9] ),
    .C(_3159_),
    .X(_3169_));
 sky130_fd_sc_hd__a21o_1 _6477_ (.A1(_1987_),
    .A2(_3157_),
    .B1(_3169_),
    .X(_0561_));
 sky130_fd_sc_hd__and3_1 _6478_ (.A(_2190_),
    .B(\immu_1.page_table[8][10] ),
    .C(_3158_),
    .X(_3170_));
 sky130_fd_sc_hd__a21o_1 _6479_ (.A1(_1989_),
    .A2(_3156_),
    .B1(_3170_),
    .X(_0562_));
 sky130_fd_sc_hd__a21bo_1 _6480_ (.A1(\inner_wb_arbiter.o_sel_sig ),
    .A2(net255),
    .B1_N(_1899_),
    .X(_3171_));
 sky130_fd_sc_hd__o211a_1 _6481_ (.A1(_1569_),
    .A2(net255),
    .B1(_3171_),
    .C1(_1911_),
    .X(_0563_));
 sky130_fd_sc_hd__nor2_8 _6482_ (.A(_1954_),
    .B(_2719_),
    .Y(_3172_));
 sky130_fd_sc_hd__mux2_1 _6483_ (.A0(\dmmu1.long_off_reg[0] ),
    .A1(_1995_),
    .S(_3172_),
    .X(_3173_));
 sky130_fd_sc_hd__clkbuf_1 _6484_ (.A(_3173_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _6485_ (.A0(\dmmu1.long_off_reg[1] ),
    .A1(_1967_),
    .S(_3172_),
    .X(_3174_));
 sky130_fd_sc_hd__clkbuf_1 _6486_ (.A(_3174_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _6487_ (.A0(\dmmu1.long_off_reg[2] ),
    .A1(_1972_),
    .S(_3172_),
    .X(_3175_));
 sky130_fd_sc_hd__clkbuf_1 _6488_ (.A(_3175_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _6489_ (.A0(\dmmu1.long_off_reg[3] ),
    .A1(_1974_),
    .S(_3172_),
    .X(_3176_));
 sky130_fd_sc_hd__clkbuf_1 _6490_ (.A(_3176_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _6491_ (.A0(\dmmu1.long_off_reg[4] ),
    .A1(_1977_),
    .S(_3172_),
    .X(_3177_));
 sky130_fd_sc_hd__clkbuf_1 _6492_ (.A(_3177_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _6493_ (.A0(\dmmu1.long_off_reg[5] ),
    .A1(_1979_),
    .S(_3172_),
    .X(_3178_));
 sky130_fd_sc_hd__clkbuf_1 _6494_ (.A(_3178_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _6495_ (.A0(\dmmu1.long_off_reg[6] ),
    .A1(_1981_),
    .S(_3172_),
    .X(_3179_));
 sky130_fd_sc_hd__clkbuf_1 _6496_ (.A(_3179_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _6497_ (.A0(\dmmu1.long_off_reg[7] ),
    .A1(_1983_),
    .S(_3172_),
    .X(_3180_));
 sky130_fd_sc_hd__clkbuf_1 _6498_ (.A(_3180_),
    .X(_0571_));
 sky130_fd_sc_hd__or3_1 _6499_ (.A(_1914_),
    .B(_1919_),
    .C(_2426_),
    .X(_3181_));
 sky130_fd_sc_hd__mux2_1 _6500_ (.A0(net96),
    .A1(\icore_sregs.c1_disable ),
    .S(_3181_),
    .X(_3182_));
 sky130_fd_sc_hd__or2_1 _6501_ (.A(net211),
    .B(_3182_),
    .X(_3183_));
 sky130_fd_sc_hd__clkbuf_1 _6502_ (.A(_3183_),
    .X(_0572_));
 sky130_fd_sc_hd__dfxtp_1 _6503_ (.CLK(clknet_leaf_60_core_clock),
    .D(_0573_),
    .Q(\immu_0.page_table[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6504_ (.CLK(clknet_leaf_59_core_clock),
    .D(_0574_),
    .Q(\immu_0.page_table[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6505_ (.CLK(clknet_leaf_62_core_clock),
    .D(_0575_),
    .Q(\immu_0.page_table[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6506_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0576_),
    .Q(\immu_0.page_table[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6507_ (.CLK(clknet_leaf_73_core_clock),
    .D(_0577_),
    .Q(\immu_0.page_table[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6508_ (.CLK(clknet_leaf_60_core_clock),
    .D(_0578_),
    .Q(\immu_0.page_table[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6509_ (.CLK(clknet_leaf_59_core_clock),
    .D(_0579_),
    .Q(\immu_0.page_table[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6510_ (.CLK(clknet_leaf_60_core_clock),
    .D(_0580_),
    .Q(\immu_0.page_table[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6511_ (.CLK(clknet_leaf_59_core_clock),
    .D(_0581_),
    .Q(\immu_0.page_table[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6512_ (.CLK(clknet_leaf_58_core_clock),
    .D(_0582_),
    .Q(\immu_0.page_table[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6513_ (.CLK(clknet_leaf_60_core_clock),
    .D(_0583_),
    .Q(\immu_0.page_table[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6514_ (.CLK(clknet_leaf_36_core_clock),
    .D(_0584_),
    .Q(\dmmu1.page_table[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6515_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0585_),
    .Q(\dmmu1.page_table[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6516_ (.CLK(clknet_leaf_36_core_clock),
    .D(_0586_),
    .Q(\dmmu1.page_table[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6517_ (.CLK(clknet_leaf_36_core_clock),
    .D(_0587_),
    .Q(\dmmu1.page_table[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6518_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0588_),
    .Q(\dmmu1.page_table[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6519_ (.CLK(clknet_leaf_36_core_clock),
    .D(_0589_),
    .Q(\dmmu1.page_table[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6520_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0590_),
    .Q(\dmmu1.page_table[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6521_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0591_),
    .Q(\dmmu1.page_table[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6522_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0592_),
    .Q(\dmmu1.page_table[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6523_ (.CLK(clknet_leaf_44_core_clock),
    .D(_0593_),
    .Q(\dmmu1.page_table[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6524_ (.CLK(clknet_leaf_31_core_clock),
    .D(_0594_),
    .Q(\dmmu1.page_table[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6525_ (.CLK(clknet_leaf_31_core_clock),
    .D(_0595_),
    .Q(\dmmu1.page_table[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6526_ (.CLK(clknet_leaf_30_core_clock),
    .D(_0596_),
    .Q(\dmmu1.page_table[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6527_ (.CLK(clknet_leaf_42_core_clock),
    .D(_0597_),
    .Q(\immu_1.page_table[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6528_ (.CLK(clknet_leaf_41_core_clock),
    .D(_0598_),
    .Q(\immu_1.page_table[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6529_ (.CLK(clknet_leaf_41_core_clock),
    .D(_0599_),
    .Q(\immu_1.page_table[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6530_ (.CLK(clknet_leaf_42_core_clock),
    .D(_0600_),
    .Q(\immu_1.page_table[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6531_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0601_),
    .Q(\immu_1.page_table[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6532_ (.CLK(clknet_leaf_46_core_clock),
    .D(_0602_),
    .Q(\immu_1.page_table[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6533_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0603_),
    .Q(\immu_1.page_table[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6534_ (.CLK(clknet_leaf_47_core_clock),
    .D(_0604_),
    .Q(\immu_1.page_table[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6535_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0605_),
    .Q(\immu_1.page_table[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6536_ (.CLK(clknet_leaf_44_core_clock),
    .D(_0606_),
    .Q(\immu_1.page_table[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6537_ (.CLK(clknet_leaf_44_core_clock),
    .D(_0607_),
    .Q(\immu_1.page_table[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6538_ (.CLK(clknet_leaf_48_core_clock),
    .D(_0608_),
    .Q(\immu_1.page_table[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6539_ (.CLK(clknet_leaf_48_core_clock),
    .D(_0609_),
    .Q(\immu_1.page_table[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6540_ (.CLK(clknet_leaf_51_core_clock),
    .D(_0610_),
    .Q(\immu_1.page_table[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6541_ (.CLK(clknet_leaf_51_core_clock),
    .D(_0611_),
    .Q(\immu_1.page_table[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6542_ (.CLK(clknet_leaf_48_core_clock),
    .D(_0612_),
    .Q(\immu_1.page_table[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6543_ (.CLK(clknet_leaf_50_core_clock),
    .D(_0613_),
    .Q(\immu_1.page_table[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6544_ (.CLK(clknet_leaf_50_core_clock),
    .D(_0614_),
    .Q(\immu_1.page_table[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6545_ (.CLK(clknet_leaf_50_core_clock),
    .D(_0615_),
    .Q(\immu_1.page_table[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6546_ (.CLK(clknet_leaf_50_core_clock),
    .D(_0616_),
    .Q(\immu_1.page_table[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6547_ (.CLK(clknet_leaf_51_core_clock),
    .D(_0617_),
    .Q(\immu_1.page_table[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6548_ (.CLK(clknet_leaf_48_core_clock),
    .D(_0618_),
    .Q(\immu_1.page_table[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6549_ (.CLK(clknet_leaf_48_core_clock),
    .D(_0619_),
    .Q(\immu_1.page_table[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6550_ (.CLK(clknet_leaf_51_core_clock),
    .D(_0620_),
    .Q(\immu_1.page_table[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6551_ (.CLK(clknet_leaf_51_core_clock),
    .D(_0621_),
    .Q(\immu_1.page_table[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6552_ (.CLK(clknet_leaf_51_core_clock),
    .D(_0622_),
    .Q(\immu_1.page_table[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6553_ (.CLK(clknet_leaf_48_core_clock),
    .D(_0623_),
    .Q(\immu_1.page_table[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6554_ (.CLK(clknet_leaf_50_core_clock),
    .D(_0624_),
    .Q(\immu_1.page_table[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6555_ (.CLK(clknet_leaf_50_core_clock),
    .D(_0625_),
    .Q(\immu_1.page_table[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6556_ (.CLK(clknet_leaf_50_core_clock),
    .D(_0626_),
    .Q(\immu_1.page_table[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6557_ (.CLK(clknet_leaf_48_core_clock),
    .D(_0627_),
    .Q(\immu_1.page_table[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6558_ (.CLK(clknet_leaf_50_core_clock),
    .D(_0628_),
    .Q(\immu_1.page_table[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6559_ (.CLK(clknet_leaf_48_core_clock),
    .D(_0629_),
    .Q(\immu_1.page_table[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6560_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0630_),
    .Q(\immu_1.page_table[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6561_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0631_),
    .Q(\immu_1.page_table[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6562_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0632_),
    .Q(\immu_1.page_table[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6563_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0633_),
    .Q(\immu_1.page_table[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6564_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0634_),
    .Q(\immu_1.page_table[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6565_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0635_),
    .Q(\immu_1.page_table[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6566_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0636_),
    .Q(\immu_1.page_table[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6567_ (.CLK(clknet_leaf_50_core_clock),
    .D(_0637_),
    .Q(\immu_1.page_table[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6568_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0638_),
    .Q(\immu_1.page_table[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6569_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0639_),
    .Q(\immu_1.page_table[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6570_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0640_),
    .Q(\immu_1.page_table[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6571_ (.CLK(clknet_leaf_46_core_clock),
    .D(_0641_),
    .Q(\immu_1.page_table[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6572_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0642_),
    .Q(\immu_1.page_table[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6573_ (.CLK(clknet_leaf_46_core_clock),
    .D(_0643_),
    .Q(\immu_1.page_table[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6574_ (.CLK(clknet_leaf_46_core_clock),
    .D(_0644_),
    .Q(\immu_1.page_table[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6575_ (.CLK(clknet_leaf_46_core_clock),
    .D(_0645_),
    .Q(\immu_1.page_table[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6576_ (.CLK(clknet_leaf_46_core_clock),
    .D(_0646_),
    .Q(\immu_1.page_table[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6577_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0647_),
    .Q(\immu_1.page_table[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6578_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0648_),
    .Q(\immu_1.page_table[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6579_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0649_),
    .Q(\immu_1.page_table[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6580_ (.CLK(clknet_leaf_49_core_clock),
    .D(_0650_),
    .Q(\immu_1.page_table[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6581_ (.CLK(clknet_leaf_46_core_clock),
    .D(_0651_),
    .Q(\immu_1.page_table[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6582_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0652_),
    .Q(\immu_1.page_table[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6583_ (.CLK(clknet_leaf_42_core_clock),
    .D(_0653_),
    .Q(\immu_1.page_table[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6584_ (.CLK(clknet_leaf_47_core_clock),
    .D(_0654_),
    .Q(\immu_1.page_table[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6585_ (.CLK(clknet_leaf_46_core_clock),
    .D(_0655_),
    .Q(\immu_1.page_table[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6586_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0656_),
    .Q(\immu_1.page_table[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6587_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0657_),
    .Q(\immu_1.page_table[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6588_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0658_),
    .Q(\immu_1.page_table[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6589_ (.CLK(clknet_leaf_44_core_clock),
    .D(_0659_),
    .Q(\immu_1.page_table[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6590_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0660_),
    .Q(\immu_1.page_table[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6591_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0661_),
    .Q(\immu_1.page_table[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6592_ (.CLK(clknet_leaf_44_core_clock),
    .D(_0662_),
    .Q(\immu_1.page_table[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6593_ (.CLK(clknet_leaf_59_core_clock),
    .D(_0663_),
    .Q(\immu_1.page_table[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6594_ (.CLK(clknet_leaf_54_core_clock),
    .D(_0664_),
    .Q(\immu_1.page_table[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6595_ (.CLK(clknet_leaf_59_core_clock),
    .D(_0665_),
    .Q(\immu_1.page_table[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6596_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0666_),
    .Q(\immu_1.page_table[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6597_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0667_),
    .Q(\immu_1.page_table[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6598_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0668_),
    .Q(\immu_1.page_table[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6599_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0669_),
    .Q(\immu_1.page_table[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6600_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0670_),
    .Q(\immu_1.page_table[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6601_ (.CLK(clknet_leaf_54_core_clock),
    .D(_0671_),
    .Q(\immu_1.page_table[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6602_ (.CLK(clknet_leaf_54_core_clock),
    .D(_0672_),
    .Q(\immu_1.page_table[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6603_ (.CLK(clknet_leaf_41_core_clock),
    .D(_0673_),
    .Q(\immu_1.page_table[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6604_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0674_),
    .Q(\immu_1.page_table[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6605_ (.CLK(clknet_leaf_54_core_clock),
    .D(_0675_),
    .Q(\immu_1.page_table[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6606_ (.CLK(clknet_leaf_62_core_clock),
    .D(_0676_),
    .Q(\immu_1.page_table[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6607_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0677_),
    .Q(\immu_1.page_table[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6608_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0678_),
    .Q(\immu_1.page_table[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6609_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0679_),
    .Q(\immu_1.page_table[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6610_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0680_),
    .Q(\immu_1.page_table[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6611_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0681_),
    .Q(\immu_1.page_table[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6612_ (.CLK(clknet_leaf_54_core_clock),
    .D(_0682_),
    .Q(\immu_1.page_table[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6613_ (.CLK(clknet_leaf_54_core_clock),
    .D(_0683_),
    .Q(\immu_1.page_table[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6614_ (.CLK(clknet_leaf_54_core_clock),
    .D(_0684_),
    .Q(\immu_1.page_table[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6615_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0685_),
    .Q(\immu_1.page_table[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6616_ (.CLK(clknet_leaf_54_core_clock),
    .D(_0686_),
    .Q(\immu_1.page_table[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6617_ (.CLK(clknet_leaf_62_core_clock),
    .D(_0687_),
    .Q(\immu_1.page_table[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6618_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0688_),
    .Q(\immu_1.page_table[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6619_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0689_),
    .Q(\immu_1.page_table[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6620_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0690_),
    .Q(\immu_1.page_table[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6621_ (.CLK(clknet_leaf_53_core_clock),
    .D(_0691_),
    .Q(\immu_1.page_table[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6622_ (.CLK(clknet_leaf_62_core_clock),
    .D(_0692_),
    .Q(\immu_1.page_table[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6623_ (.CLK(clknet_leaf_54_core_clock),
    .D(_0693_),
    .Q(\immu_1.page_table[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6624_ (.CLK(clknet_leaf_54_core_clock),
    .D(_0694_),
    .Q(\immu_1.page_table[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6625_ (.CLK(clknet_leaf_54_core_clock),
    .D(_0695_),
    .Q(\immu_1.page_table[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6626_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0696_),
    .Q(\immu_1.page_table[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6627_ (.CLK(clknet_leaf_41_core_clock),
    .D(_0697_),
    .Q(\immu_1.page_table[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6628_ (.CLK(clknet_leaf_55_core_clock),
    .D(_0698_),
    .Q(\immu_1.page_table[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6629_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0699_),
    .Q(\immu_1.page_table[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6630_ (.CLK(clknet_leaf_55_core_clock),
    .D(_0700_),
    .Q(\immu_1.page_table[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6631_ (.CLK(clknet_leaf_55_core_clock),
    .D(_0701_),
    .Q(\immu_1.page_table[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6632_ (.CLK(clknet_leaf_41_core_clock),
    .D(_0702_),
    .Q(\immu_1.page_table[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6633_ (.CLK(clknet_leaf_40_core_clock),
    .D(_0703_),
    .Q(\immu_1.page_table[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6634_ (.CLK(clknet_leaf_40_core_clock),
    .D(_0704_),
    .Q(\immu_1.page_table[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6635_ (.CLK(clknet_leaf_40_core_clock),
    .D(_0705_),
    .Q(\immu_1.page_table[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6636_ (.CLK(clknet_leaf_40_core_clock),
    .D(_0706_),
    .Q(\immu_1.page_table[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6637_ (.CLK(clknet_leaf_57_core_clock),
    .D(_0707_),
    .Q(\immu_1.page_table[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6638_ (.CLK(clknet_leaf_42_core_clock),
    .D(_0708_),
    .Q(\immu_1.page_table[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6639_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0709_),
    .Q(\immu_1.page_table[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6640_ (.CLK(clknet_leaf_57_core_clock),
    .D(_0710_),
    .Q(\immu_1.page_table[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6641_ (.CLK(clknet_leaf_38_core_clock),
    .D(_0711_),
    .Q(\immu_1.page_table[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6642_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0712_),
    .Q(\immu_1.page_table[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6643_ (.CLK(clknet_leaf_39_core_clock),
    .D(_0713_),
    .Q(\immu_1.page_table[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6644_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0714_),
    .Q(\immu_1.page_table[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6645_ (.CLK(clknet_leaf_40_core_clock),
    .D(_0715_),
    .Q(\immu_1.page_table[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6646_ (.CLK(clknet_leaf_42_core_clock),
    .D(_0716_),
    .Q(\immu_1.page_table[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6647_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0717_),
    .Q(\immu_1.page_table[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6648_ (.CLK(clknet_leaf_38_core_clock),
    .D(_0718_),
    .Q(\immu_1.page_table[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6649_ (.CLK(clknet_leaf_40_core_clock),
    .D(_0719_),
    .Q(\immu_1.page_table[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6650_ (.CLK(clknet_leaf_39_core_clock),
    .D(_0720_),
    .Q(\immu_1.page_table[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6651_ (.CLK(clknet_leaf_38_core_clock),
    .D(_0721_),
    .Q(\immu_1.page_table[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6652_ (.CLK(clknet_leaf_38_core_clock),
    .D(_0722_),
    .Q(\immu_1.page_table[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6653_ (.CLK(clknet_leaf_39_core_clock),
    .D(_0723_),
    .Q(\immu_1.page_table[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6654_ (.CLK(clknet_leaf_40_core_clock),
    .D(_0724_),
    .Q(\immu_1.page_table[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6655_ (.CLK(clknet_leaf_39_core_clock),
    .D(_0725_),
    .Q(\immu_1.page_table[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6656_ (.CLK(clknet_leaf_40_core_clock),
    .D(_0726_),
    .Q(\immu_1.page_table[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6657_ (.CLK(clknet_leaf_42_core_clock),
    .D(_0727_),
    .Q(\immu_1.page_table[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6658_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0728_),
    .Q(\immu_1.page_table[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6659_ (.CLK(clknet_leaf_8_core_clock),
    .D(_0729_),
    .Q(\dmmu0.page_table[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6660_ (.CLK(clknet_leaf_7_core_clock),
    .D(_0730_),
    .Q(\dmmu0.page_table[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6661_ (.CLK(clknet_leaf_80_core_clock),
    .D(_0731_),
    .Q(\dmmu0.page_table[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6662_ (.CLK(clknet_leaf_80_core_clock),
    .D(_0732_),
    .Q(\dmmu0.page_table[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6663_ (.CLK(clknet_leaf_9_core_clock),
    .D(_0733_),
    .Q(\dmmu0.page_table[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6664_ (.CLK(clknet_leaf_8_core_clock),
    .D(_0734_),
    .Q(\dmmu0.page_table[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6665_ (.CLK(clknet_leaf_9_core_clock),
    .D(_0735_),
    .Q(\dmmu0.page_table[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6666_ (.CLK(clknet_leaf_8_core_clock),
    .D(_0736_),
    .Q(\dmmu0.page_table[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6667_ (.CLK(clknet_leaf_9_core_clock),
    .D(_0737_),
    .Q(\dmmu0.page_table[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6668_ (.CLK(clknet_leaf_5_core_clock),
    .D(_0738_),
    .Q(\dmmu0.page_table[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6669_ (.CLK(clknet_leaf_3_core_clock),
    .D(_0739_),
    .Q(\dmmu0.page_table[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6670_ (.CLK(clknet_leaf_2_core_clock),
    .D(_0740_),
    .Q(\dmmu0.page_table[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6671_ (.CLK(clknet_leaf_4_core_clock),
    .D(_0741_),
    .Q(\dmmu0.page_table[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6672_ (.CLK(clknet_leaf_58_core_clock),
    .D(_0742_),
    .Q(\immu_1.page_table[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6673_ (.CLK(clknet_leaf_58_core_clock),
    .D(_0743_),
    .Q(\immu_1.page_table[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6674_ (.CLK(clknet_leaf_58_core_clock),
    .D(_0744_),
    .Q(\immu_1.page_table[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6675_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0745_),
    .Q(\immu_1.page_table[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6676_ (.CLK(clknet_leaf_55_core_clock),
    .D(_0746_),
    .Q(\immu_1.page_table[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6677_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0747_),
    .Q(\immu_1.page_table[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6678_ (.CLK(clknet_leaf_55_core_clock),
    .D(_0748_),
    .Q(\immu_1.page_table[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6679_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0749_),
    .Q(\immu_1.page_table[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6680_ (.CLK(clknet_leaf_54_core_clock),
    .D(_0750_),
    .Q(\immu_1.page_table[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6681_ (.CLK(clknet_leaf_41_core_clock),
    .D(_0751_),
    .Q(\immu_1.page_table[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6682_ (.CLK(clknet_leaf_41_core_clock),
    .D(_0752_),
    .Q(\immu_1.page_table[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6683_ (.CLK(clknet_leaf_40_core_clock),
    .D(_0753_),
    .Q(\immu_1.page_table[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6684_ (.CLK(clknet_leaf_42_core_clock),
    .D(_0754_),
    .Q(\immu_1.page_table[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6685_ (.CLK(clknet_leaf_57_core_clock),
    .D(_0755_),
    .Q(\immu_1.page_table[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6686_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0756_),
    .Q(\immu_1.page_table[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6687_ (.CLK(clknet_leaf_39_core_clock),
    .D(_0757_),
    .Q(\immu_1.page_table[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6688_ (.CLK(clknet_leaf_56_core_clock),
    .D(_0758_),
    .Q(\immu_1.page_table[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6689_ (.CLK(clknet_leaf_39_core_clock),
    .D(_0759_),
    .Q(\immu_1.page_table[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6690_ (.CLK(clknet_leaf_58_core_clock),
    .D(_0760_),
    .Q(\immu_1.page_table[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6691_ (.CLK(clknet_leaf_39_core_clock),
    .D(_0761_),
    .Q(\immu_1.page_table[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6692_ (.CLK(clknet_leaf_42_core_clock),
    .D(_0762_),
    .Q(\immu_1.page_table[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6693_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0763_),
    .Q(\immu_1.page_table[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6694_ (.CLK(clknet_leaf_41_core_clock),
    .D(_0764_),
    .Q(\immu_1.page_table[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6695_ (.CLK(clknet_leaf_42_core_clock),
    .D(_0765_),
    .Q(\immu_1.page_table[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6696_ (.CLK(clknet_leaf_41_core_clock),
    .D(_0766_),
    .Q(\immu_1.page_table[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6697_ (.CLK(clknet_leaf_42_core_clock),
    .D(_0767_),
    .Q(\immu_1.page_table[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6698_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0768_),
    .Q(\immu_1.page_table[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6699_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0769_),
    .Q(\immu_1.page_table[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6700_ (.CLK(clknet_leaf_42_core_clock),
    .D(_0770_),
    .Q(\immu_1.page_table[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6701_ (.CLK(clknet_leaf_42_core_clock),
    .D(_0771_),
    .Q(\immu_1.page_table[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6702_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0772_),
    .Q(\immu_1.page_table[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6703_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0773_),
    .Q(\immu_1.page_table[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6704_ (.CLK(clknet_leaf_45_core_clock),
    .D(_0774_),
    .Q(\immu_1.page_table[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6705_ (.CLK(clknet_leaf_62_core_clock),
    .D(_0775_),
    .Q(\immu_0.page_table[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6706_ (.CLK(clknet_leaf_61_core_clock),
    .D(_0776_),
    .Q(\immu_0.page_table[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6707_ (.CLK(clknet_leaf_62_core_clock),
    .D(_0777_),
    .Q(\immu_0.page_table[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6708_ (.CLK(clknet_leaf_61_core_clock),
    .D(_0778_),
    .Q(\immu_0.page_table[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6709_ (.CLK(clknet_leaf_63_core_clock),
    .D(_0779_),
    .Q(\immu_0.page_table[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6710_ (.CLK(clknet_leaf_63_core_clock),
    .D(_0780_),
    .Q(\immu_0.page_table[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6711_ (.CLK(clknet_leaf_61_core_clock),
    .D(_0781_),
    .Q(\immu_0.page_table[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6712_ (.CLK(clknet_leaf_63_core_clock),
    .D(_0782_),
    .Q(\immu_0.page_table[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6713_ (.CLK(clknet_leaf_61_core_clock),
    .D(_0783_),
    .Q(\immu_0.page_table[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6714_ (.CLK(clknet_leaf_62_core_clock),
    .D(_0784_),
    .Q(\immu_0.page_table[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6715_ (.CLK(clknet_leaf_61_core_clock),
    .D(_0785_),
    .Q(\immu_0.page_table[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6716_ (.CLK(clknet_leaf_62_core_clock),
    .D(_0786_),
    .Q(\immu_0.page_table[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6717_ (.CLK(clknet_leaf_63_core_clock),
    .D(_0787_),
    .Q(\immu_0.page_table[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6718_ (.CLK(clknet_leaf_62_core_clock),
    .D(_0788_),
    .Q(\immu_0.page_table[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6719_ (.CLK(clknet_leaf_63_core_clock),
    .D(_0789_),
    .Q(\immu_0.page_table[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6720_ (.CLK(clknet_leaf_63_core_clock),
    .D(_0790_),
    .Q(\immu_0.page_table[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6721_ (.CLK(clknet_leaf_63_core_clock),
    .D(_0791_),
    .Q(\immu_0.page_table[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6722_ (.CLK(clknet_leaf_67_core_clock),
    .D(_0792_),
    .Q(\immu_0.page_table[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6723_ (.CLK(clknet_leaf_63_core_clock),
    .D(_0793_),
    .Q(\immu_0.page_table[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6724_ (.CLK(clknet_leaf_61_core_clock),
    .D(_0794_),
    .Q(\immu_0.page_table[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6725_ (.CLK(clknet_leaf_62_core_clock),
    .D(_0795_),
    .Q(\immu_0.page_table[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6726_ (.CLK(clknet_leaf_61_core_clock),
    .D(_0796_),
    .Q(\immu_0.page_table[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6727_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0797_),
    .Q(\immu_0.page_table[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6728_ (.CLK(clknet_3_2_0_core_clock),
    .D(_0798_),
    .Q(\immu_0.page_table[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6729_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0799_),
    .Q(\immu_0.page_table[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6730_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0800_),
    .Q(\immu_0.page_table[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6731_ (.CLK(clknet_leaf_67_core_clock),
    .D(_0801_),
    .Q(\immu_0.page_table[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6732_ (.CLK(clknet_leaf_63_core_clock),
    .D(_0802_),
    .Q(\immu_0.page_table[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6733_ (.CLK(clknet_leaf_63_core_clock),
    .D(_0803_),
    .Q(\immu_0.page_table[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6734_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0804_),
    .Q(\immu_0.page_table[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6735_ (.CLK(clknet_leaf_67_core_clock),
    .D(_0805_),
    .Q(\immu_0.page_table[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6736_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0806_),
    .Q(\immu_0.page_table[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6737_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0807_),
    .Q(\immu_0.page_table[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6738_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0808_),
    .Q(\immu_0.page_table[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6739_ (.CLK(clknet_leaf_67_core_clock),
    .D(_0000_),
    .Q(\immu_0.page_table[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6740_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0001_),
    .Q(\immu_0.page_table[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6741_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0002_),
    .Q(\immu_0.page_table[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6742_ (.CLK(clknet_leaf_67_core_clock),
    .D(_0003_),
    .Q(\immu_0.page_table[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6743_ (.CLK(clknet_leaf_67_core_clock),
    .D(_0004_),
    .Q(\immu_0.page_table[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6744_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0005_),
    .Q(\immu_0.page_table[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6745_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0006_),
    .Q(\immu_0.page_table[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6746_ (.CLK(clknet_leaf_67_core_clock),
    .D(_0007_),
    .Q(\immu_0.page_table[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6747_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0008_),
    .Q(\immu_0.page_table[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6748_ (.CLK(clknet_leaf_67_core_clock),
    .D(_0009_),
    .Q(\immu_0.page_table[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6749_ (.CLK(clknet_leaf_87_core_clock),
    .D(_0010_),
    .Q(\dmmu0.page_table[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6750_ (.CLK(clknet_leaf_89_core_clock),
    .D(_0011_),
    .Q(\dmmu0.page_table[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6751_ (.CLK(clknet_leaf_88_core_clock),
    .D(_0012_),
    .Q(\dmmu0.page_table[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6752_ (.CLK(clknet_leaf_86_core_clock),
    .D(_0013_),
    .Q(\dmmu0.page_table[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6753_ (.CLK(clknet_leaf_88_core_clock),
    .D(_0014_),
    .Q(\dmmu0.page_table[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6754_ (.CLK(clknet_leaf_89_core_clock),
    .D(_0015_),
    .Q(\dmmu0.page_table[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6755_ (.CLK(clknet_leaf_89_core_clock),
    .D(_0016_),
    .Q(\dmmu0.page_table[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6756_ (.CLK(clknet_leaf_90_core_clock),
    .D(_0017_),
    .Q(\dmmu0.page_table[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6757_ (.CLK(clknet_leaf_90_core_clock),
    .D(_0018_),
    .Q(\dmmu0.page_table[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6758_ (.CLK(clknet_leaf_89_core_clock),
    .D(_0019_),
    .Q(\dmmu0.page_table[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6759_ (.CLK(clknet_leaf_93_core_clock),
    .D(_0020_),
    .Q(\dmmu0.page_table[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6760_ (.CLK(clknet_leaf_0_core_clock),
    .D(_0021_),
    .Q(\dmmu0.page_table[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6761_ (.CLK(clknet_leaf_93_core_clock),
    .D(_0022_),
    .Q(\dmmu0.page_table[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6762_ (.CLK(clknet_leaf_87_core_clock),
    .D(_0023_),
    .Q(\dmmu0.page_table[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6763_ (.CLK(clknet_leaf_86_core_clock),
    .D(_0024_),
    .Q(\dmmu0.page_table[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6764_ (.CLK(clknet_leaf_87_core_clock),
    .D(_0025_),
    .Q(\dmmu0.page_table[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6765_ (.CLK(clknet_leaf_85_core_clock),
    .D(_0026_),
    .Q(\dmmu0.page_table[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6766_ (.CLK(clknet_leaf_87_core_clock),
    .D(_0027_),
    .Q(\dmmu0.page_table[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6767_ (.CLK(clknet_leaf_89_core_clock),
    .D(_0028_),
    .Q(\dmmu0.page_table[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6768_ (.CLK(clknet_leaf_86_core_clock),
    .D(_0029_),
    .Q(\dmmu0.page_table[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6769_ (.CLK(clknet_leaf_90_core_clock),
    .D(_0030_),
    .Q(\dmmu0.page_table[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6770_ (.CLK(clknet_leaf_90_core_clock),
    .D(_0031_),
    .Q(\dmmu0.page_table[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6771_ (.CLK(clknet_leaf_89_core_clock),
    .D(_0032_),
    .Q(\dmmu0.page_table[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6772_ (.CLK(clknet_leaf_91_core_clock),
    .D(_0033_),
    .Q(\dmmu0.page_table[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6773_ (.CLK(clknet_leaf_91_core_clock),
    .D(_0034_),
    .Q(\dmmu0.page_table[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6774_ (.CLK(clknet_leaf_91_core_clock),
    .D(_0035_),
    .Q(\dmmu0.page_table[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6775_ (.CLK(clknet_leaf_81_core_clock),
    .D(_0036_),
    .Q(\dmmu0.page_table[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6776_ (.CLK(clknet_leaf_85_core_clock),
    .D(_0037_),
    .Q(\dmmu0.page_table[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6777_ (.CLK(clknet_leaf_81_core_clock),
    .D(_0038_),
    .Q(\dmmu0.page_table[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6778_ (.CLK(clknet_leaf_85_core_clock),
    .D(_0039_),
    .Q(\dmmu0.page_table[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6779_ (.CLK(clknet_leaf_87_core_clock),
    .D(_0040_),
    .Q(\dmmu0.page_table[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6780_ (.CLK(clknet_leaf_89_core_clock),
    .D(_0041_),
    .Q(\dmmu0.page_table[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6781_ (.CLK(clknet_leaf_86_core_clock),
    .D(_0042_),
    .Q(\dmmu0.page_table[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6782_ (.CLK(clknet_leaf_89_core_clock),
    .D(_0043_),
    .Q(\dmmu0.page_table[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6783_ (.CLK(clknet_leaf_90_core_clock),
    .D(_0044_),
    .Q(\dmmu0.page_table[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6784_ (.CLK(clknet_leaf_89_core_clock),
    .D(_0045_),
    .Q(\dmmu0.page_table[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6785_ (.CLK(clknet_leaf_0_core_clock),
    .D(_0046_),
    .Q(\dmmu0.page_table[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6786_ (.CLK(clknet_leaf_0_core_clock),
    .D(_0047_),
    .Q(\dmmu0.page_table[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6787_ (.CLK(clknet_leaf_0_core_clock),
    .D(_0048_),
    .Q(\dmmu0.page_table[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 _6788_ (.CLK(clknet_leaf_2_core_clock),
    .D(_0049_),
    .Q(net407));
 sky130_fd_sc_hd__dfxtp_2 _6789_ (.CLK(clknet_leaf_3_core_clock),
    .D(_0050_),
    .Q(net408));
 sky130_fd_sc_hd__dfxtp_1 _6790_ (.CLK(clknet_leaf_80_core_clock),
    .D(_0051_),
    .Q(\dmmu0.page_table[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6791_ (.CLK(clknet_leaf_80_core_clock),
    .D(_0052_),
    .Q(\dmmu0.page_table[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6792_ (.CLK(clknet_leaf_80_core_clock),
    .D(_0053_),
    .Q(\dmmu0.page_table[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6793_ (.CLK(clknet_leaf_80_core_clock),
    .D(_0054_),
    .Q(\dmmu0.page_table[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6794_ (.CLK(clknet_leaf_10_core_clock),
    .D(_0055_),
    .Q(\dmmu0.page_table[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6795_ (.CLK(clknet_leaf_80_core_clock),
    .D(_0056_),
    .Q(\dmmu0.page_table[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6796_ (.CLK(clknet_leaf_10_core_clock),
    .D(_0057_),
    .Q(\dmmu0.page_table[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6797_ (.CLK(clknet_leaf_10_core_clock),
    .D(_0058_),
    .Q(\dmmu0.page_table[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6798_ (.CLK(clknet_leaf_10_core_clock),
    .D(_0059_),
    .Q(\dmmu0.page_table[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6799_ (.CLK(clknet_leaf_8_core_clock),
    .D(_0060_),
    .Q(\dmmu0.page_table[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6800_ (.CLK(clknet_leaf_6_core_clock),
    .D(_0061_),
    .Q(\dmmu0.page_table[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6801_ (.CLK(clknet_leaf_6_core_clock),
    .D(_0062_),
    .Q(\dmmu0.page_table[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6802_ (.CLK(clknet_leaf_6_core_clock),
    .D(_0063_),
    .Q(\dmmu0.page_table[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6803_ (.CLK(clknet_leaf_81_core_clock),
    .D(_0064_),
    .Q(\dmmu0.page_table[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6804_ (.CLK(clknet_leaf_84_core_clock),
    .D(_0065_),
    .Q(\dmmu0.page_table[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6805_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0066_),
    .Q(\dmmu0.page_table[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6806_ (.CLK(clknet_leaf_84_core_clock),
    .D(_0067_),
    .Q(\dmmu0.page_table[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6807_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0068_),
    .Q(\dmmu0.page_table[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6808_ (.CLK(clknet_leaf_85_core_clock),
    .D(_0069_),
    .Q(\dmmu0.page_table[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6809_ (.CLK(clknet_leaf_86_core_clock),
    .D(_0070_),
    .Q(\dmmu0.page_table[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6810_ (.CLK(clknet_leaf_87_core_clock),
    .D(_0071_),
    .Q(\dmmu0.page_table[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6811_ (.CLK(clknet_leaf_85_core_clock),
    .D(_0072_),
    .Q(\dmmu0.page_table[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6812_ (.CLK(clknet_leaf_87_core_clock),
    .D(_0073_),
    .Q(\dmmu0.page_table[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6813_ (.CLK(clknet_leaf_1_core_clock),
    .D(_0074_),
    .Q(\dmmu0.page_table[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6814_ (.CLK(clknet_leaf_88_core_clock),
    .D(_0075_),
    .Q(\dmmu0.page_table[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6815_ (.CLK(clknet_leaf_0_core_clock),
    .D(_0076_),
    .Q(\dmmu0.page_table[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6816_ (.CLK(clknet_leaf_60_core_clock),
    .D(_0077_),
    .Q(\immu_0.page_table[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6817_ (.CLK(clknet_leaf_59_core_clock),
    .D(_0078_),
    .Q(\immu_0.page_table[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6818_ (.CLK(clknet_leaf_59_core_clock),
    .D(_0079_),
    .Q(\immu_0.page_table[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6819_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0080_),
    .Q(\immu_0.page_table[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6820_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0081_),
    .Q(\immu_0.page_table[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6821_ (.CLK(clknet_leaf_61_core_clock),
    .D(_0082_),
    .Q(\immu_0.page_table[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6822_ (.CLK(clknet_leaf_59_core_clock),
    .D(_0083_),
    .Q(\immu_0.page_table[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6823_ (.CLK(clknet_leaf_74_core_clock),
    .D(_0084_),
    .Q(\immu_0.page_table[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6824_ (.CLK(clknet_leaf_59_core_clock),
    .D(_0085_),
    .Q(\immu_0.page_table[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6825_ (.CLK(clknet_leaf_59_core_clock),
    .D(_0086_),
    .Q(\immu_0.page_table[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6826_ (.CLK(clknet_leaf_60_core_clock),
    .D(_0087_),
    .Q(\immu_0.page_table[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6827_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0088_),
    .Q(\immu_0.page_table[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6828_ (.CLK(clknet_leaf_73_core_clock),
    .D(_0089_),
    .Q(\immu_0.page_table[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6829_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0090_),
    .Q(\immu_0.page_table[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6830_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0091_),
    .Q(\immu_0.page_table[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6831_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0092_),
    .Q(\immu_0.page_table[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6832_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0093_),
    .Q(\immu_0.page_table[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6833_ (.CLK(clknet_leaf_66_core_clock),
    .D(_0094_),
    .Q(\immu_0.page_table[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6834_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0095_),
    .Q(\immu_0.page_table[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6835_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0096_),
    .Q(\immu_0.page_table[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6836_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0097_),
    .Q(\immu_0.page_table[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6837_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0098_),
    .Q(\immu_0.page_table[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6838_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0099_),
    .Q(\immu_0.page_table[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6839_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0100_),
    .Q(\immu_0.page_table[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6840_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0101_),
    .Q(\immu_0.page_table[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6841_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0102_),
    .Q(\immu_0.page_table[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6842_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0103_),
    .Q(\immu_0.page_table[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6843_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0104_),
    .Q(\immu_0.page_table[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6844_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0105_),
    .Q(\immu_0.page_table[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6845_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0106_),
    .Q(\immu_0.page_table[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6846_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0107_),
    .Q(\immu_0.page_table[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6847_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0108_),
    .Q(\immu_0.page_table[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6848_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0109_),
    .Q(\immu_0.page_table[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6849_ (.CLK(clknet_leaf_73_core_clock),
    .D(_0110_),
    .Q(\immu_0.page_table[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6850_ (.CLK(clknet_leaf_70_core_clock),
    .D(_0111_),
    .Q(\immu_0.page_table[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6851_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0112_),
    .Q(\immu_0.page_table[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6852_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0113_),
    .Q(\immu_0.page_table[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6853_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0114_),
    .Q(\immu_0.page_table[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6854_ (.CLK(clknet_leaf_70_core_clock),
    .D(_0115_),
    .Q(\immu_0.page_table[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6855_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0116_),
    .Q(\immu_0.page_table[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6856_ (.CLK(clknet_leaf_68_core_clock),
    .D(_0117_),
    .Q(\immu_0.page_table[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6857_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0118_),
    .Q(\immu_0.page_table[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6858_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0119_),
    .Q(\immu_0.page_table[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6859_ (.CLK(clknet_leaf_72_core_clock),
    .D(_0120_),
    .Q(\immu_0.page_table[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6860_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0121_),
    .Q(\immu_0.page_table[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6861_ (.CLK(clknet_leaf_70_core_clock),
    .D(_0122_),
    .Q(\immu_0.page_table[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6862_ (.CLK(clknet_leaf_70_core_clock),
    .D(_0123_),
    .Q(\immu_0.page_table[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6863_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0124_),
    .Q(\immu_0.page_table[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6864_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0125_),
    .Q(\immu_0.page_table[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6865_ (.CLK(clknet_leaf_70_core_clock),
    .D(_0126_),
    .Q(\immu_0.page_table[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6866_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0127_),
    .Q(\immu_0.page_table[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6867_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0128_),
    .Q(\immu_0.page_table[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6868_ (.CLK(clknet_leaf_73_core_clock),
    .D(_0129_),
    .Q(\immu_0.page_table[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6869_ (.CLK(clknet_leaf_69_core_clock),
    .D(_0130_),
    .Q(\immu_0.page_table[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6870_ (.CLK(clknet_leaf_72_core_clock),
    .D(_0131_),
    .Q(\immu_0.page_table[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6871_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0132_),
    .Q(\immu_0.page_table[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6872_ (.CLK(clknet_leaf_70_core_clock),
    .D(_0133_),
    .Q(\immu_0.page_table[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6873_ (.CLK(clknet_leaf_70_core_clock),
    .D(_0134_),
    .Q(\immu_0.page_table[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6874_ (.CLK(clknet_leaf_70_core_clock),
    .D(_0135_),
    .Q(\immu_0.page_table[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6875_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0136_),
    .Q(\immu_0.page_table[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6876_ (.CLK(clknet_leaf_70_core_clock),
    .D(_0137_),
    .Q(\immu_0.page_table[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6877_ (.CLK(clknet_leaf_70_core_clock),
    .D(_0138_),
    .Q(\immu_0.page_table[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6878_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0139_),
    .Q(\immu_0.page_table[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6879_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0140_),
    .Q(\immu_0.page_table[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6880_ (.CLK(clknet_leaf_70_core_clock),
    .D(_0141_),
    .Q(\immu_0.page_table[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6881_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0142_),
    .Q(\immu_0.page_table[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6882_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0143_),
    .Q(\immu_0.page_table[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6883_ (.CLK(clknet_leaf_84_core_clock),
    .D(_0144_),
    .Q(\immu_0.page_table[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6884_ (.CLK(clknet_leaf_84_core_clock),
    .D(_0145_),
    .Q(\immu_0.page_table[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6885_ (.CLK(clknet_leaf_84_core_clock),
    .D(_0146_),
    .Q(\immu_0.page_table[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6886_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0147_),
    .Q(\immu_0.page_table[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6887_ (.CLK(clknet_leaf_84_core_clock),
    .D(_0148_),
    .Q(\immu_0.page_table[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6888_ (.CLK(clknet_leaf_83_core_clock),
    .D(_0149_),
    .Q(\immu_0.page_table[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6889_ (.CLK(clknet_leaf_83_core_clock),
    .D(_0150_),
    .Q(\immu_0.page_table[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6890_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0151_),
    .Q(\immu_0.page_table[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6891_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0152_),
    .Q(\immu_0.page_table[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6892_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0153_),
    .Q(\immu_0.page_table[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6893_ (.CLK(clknet_leaf_76_core_clock),
    .D(_0154_),
    .Q(\immu_0.page_table[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6894_ (.CLK(clknet_leaf_72_core_clock),
    .D(_0155_),
    .Q(\immu_0.page_table[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6895_ (.CLK(clknet_leaf_71_core_clock),
    .D(_0156_),
    .Q(\immu_0.page_table[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6896_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0157_),
    .Q(\immu_0.page_table[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6897_ (.CLK(clknet_leaf_75_core_clock),
    .D(_0158_),
    .Q(\immu_0.page_table[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6898_ (.CLK(clknet_leaf_76_core_clock),
    .D(_0159_),
    .Q(\immu_0.page_table[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6899_ (.CLK(clknet_leaf_76_core_clock),
    .D(_0160_),
    .Q(\immu_0.page_table[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6900_ (.CLK(clknet_leaf_75_core_clock),
    .D(_0161_),
    .Q(\immu_0.page_table[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6901_ (.CLK(clknet_leaf_72_core_clock),
    .D(_0162_),
    .Q(\immu_0.page_table[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6902_ (.CLK(clknet_leaf_79_core_clock),
    .D(_0163_),
    .Q(\immu_0.page_table[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6903_ (.CLK(clknet_leaf_76_core_clock),
    .D(_0164_),
    .Q(\immu_0.page_table[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6904_ (.CLK(clknet_leaf_79_core_clock),
    .D(_0165_),
    .Q(\immu_0.page_table[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6905_ (.CLK(clknet_leaf_72_core_clock),
    .D(_0166_),
    .Q(\immu_0.page_table[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6906_ (.CLK(clknet_leaf_72_core_clock),
    .D(_0167_),
    .Q(\immu_0.page_table[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6907_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0168_),
    .Q(\immu_0.page_table[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6908_ (.CLK(clknet_leaf_75_core_clock),
    .D(_0169_),
    .Q(\immu_0.page_table[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6909_ (.CLK(clknet_leaf_76_core_clock),
    .D(_0170_),
    .Q(\immu_0.page_table[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6910_ (.CLK(clknet_leaf_76_core_clock),
    .D(_0171_),
    .Q(\immu_0.page_table[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6911_ (.CLK(clknet_leaf_76_core_clock),
    .D(_0172_),
    .Q(\immu_0.page_table[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6912_ (.CLK(clknet_leaf_72_core_clock),
    .D(_0173_),
    .Q(\immu_0.page_table[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6913_ (.CLK(clknet_leaf_79_core_clock),
    .D(_0174_),
    .Q(\immu_0.page_table[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6914_ (.CLK(clknet_leaf_79_core_clock),
    .D(_0175_),
    .Q(\immu_0.page_table[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6915_ (.CLK(clknet_leaf_76_core_clock),
    .D(_0176_),
    .Q(\immu_0.page_table[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6916_ (.CLK(clknet_leaf_74_core_clock),
    .D(_0177_),
    .Q(\immu_0.page_table[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6917_ (.CLK(clknet_leaf_58_core_clock),
    .D(_0178_),
    .Q(\immu_0.page_table[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6918_ (.CLK(clknet_leaf_75_core_clock),
    .D(_0179_),
    .Q(\immu_0.page_table[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6919_ (.CLK(clknet_leaf_75_core_clock),
    .D(_0180_),
    .Q(\immu_0.page_table[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6920_ (.CLK(clknet_leaf_76_core_clock),
    .D(_0181_),
    .Q(\immu_0.page_table[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6921_ (.CLK(clknet_leaf_57_core_clock),
    .D(_0182_),
    .Q(\immu_0.page_table[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6922_ (.CLK(clknet_leaf_77_core_clock),
    .D(_0183_),
    .Q(\immu_0.page_table[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6923_ (.CLK(clknet_leaf_75_core_clock),
    .D(_0184_),
    .Q(\immu_0.page_table[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6924_ (.CLK(clknet_leaf_58_core_clock),
    .D(_0185_),
    .Q(\immu_0.page_table[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6925_ (.CLK(clknet_leaf_77_core_clock),
    .D(_0186_),
    .Q(\immu_0.page_table[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6926_ (.CLK(clknet_leaf_76_core_clock),
    .D(_0187_),
    .Q(\immu_0.page_table[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6927_ (.CLK(clknet_leaf_60_core_clock),
    .D(_0188_),
    .Q(\immu_0.page_table[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6928_ (.CLK(clknet_leaf_58_core_clock),
    .D(_0189_),
    .Q(\immu_0.page_table[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6929_ (.CLK(clknet_leaf_77_core_clock),
    .D(_0190_),
    .Q(\immu_0.page_table[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6930_ (.CLK(clknet_leaf_77_core_clock),
    .D(_0191_),
    .Q(\immu_0.page_table[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6931_ (.CLK(clknet_leaf_77_core_clock),
    .D(_0192_),
    .Q(\immu_0.page_table[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6932_ (.CLK(clknet_leaf_57_core_clock),
    .D(_0193_),
    .Q(\immu_0.page_table[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6933_ (.CLK(clknet_leaf_57_core_clock),
    .D(_0194_),
    .Q(\immu_0.page_table[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6934_ (.CLK(clknet_leaf_75_core_clock),
    .D(_0195_),
    .Q(\immu_0.page_table[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6935_ (.CLK(clknet_leaf_58_core_clock),
    .D(_0196_),
    .Q(\immu_0.page_table[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6936_ (.CLK(clknet_leaf_77_core_clock),
    .D(_0197_),
    .Q(\immu_0.page_table[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6937_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0198_),
    .Q(\dmmu0.page_table[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6938_ (.CLK(clknet_leaf_84_core_clock),
    .D(_0199_),
    .Q(\dmmu0.page_table[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6939_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0200_),
    .Q(\dmmu0.page_table[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6940_ (.CLK(clknet_leaf_84_core_clock),
    .D(_0201_),
    .Q(\dmmu0.page_table[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6941_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0202_),
    .Q(\dmmu0.page_table[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6942_ (.CLK(clknet_leaf_85_core_clock),
    .D(_0203_),
    .Q(\dmmu0.page_table[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6943_ (.CLK(clknet_leaf_85_core_clock),
    .D(_0204_),
    .Q(\dmmu0.page_table[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6944_ (.CLK(clknet_leaf_83_core_clock),
    .D(_0205_),
    .Q(\dmmu0.page_table[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6945_ (.CLK(clknet_leaf_85_core_clock),
    .D(_0206_),
    .Q(\dmmu0.page_table[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6946_ (.CLK(clknet_leaf_81_core_clock),
    .D(_0207_),
    .Q(\dmmu0.page_table[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6947_ (.CLK(clknet_leaf_1_core_clock),
    .D(_0208_),
    .Q(\dmmu0.page_table[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6948_ (.CLK(clknet_leaf_81_core_clock),
    .D(_0209_),
    .Q(\dmmu0.page_table[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6949_ (.CLK(clknet_leaf_7_core_clock),
    .D(_0210_),
    .Q(\dmmu0.page_table[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6950_ (.CLK(clknet_leaf_81_core_clock),
    .D(_0211_),
    .Q(\dmmu0.page_table[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6951_ (.CLK(clknet_leaf_84_core_clock),
    .D(_0212_),
    .Q(\dmmu0.page_table[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6952_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0213_),
    .Q(\dmmu0.page_table[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6953_ (.CLK(clknet_leaf_84_core_clock),
    .D(_0214_),
    .Q(\dmmu0.page_table[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6954_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0215_),
    .Q(\dmmu0.page_table[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6955_ (.CLK(clknet_leaf_85_core_clock),
    .D(_0216_),
    .Q(\dmmu0.page_table[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6956_ (.CLK(clknet_leaf_85_core_clock),
    .D(_0217_),
    .Q(\dmmu0.page_table[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6957_ (.CLK(clknet_leaf_81_core_clock),
    .D(_0218_),
    .Q(\dmmu0.page_table[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6958_ (.CLK(clknet_leaf_85_core_clock),
    .D(_0219_),
    .Q(\dmmu0.page_table[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6959_ (.CLK(clknet_leaf_87_core_clock),
    .D(_0220_),
    .Q(\dmmu0.page_table[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6960_ (.CLK(clknet_leaf_88_core_clock),
    .D(_0221_),
    .Q(\dmmu0.page_table[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6961_ (.CLK(clknet_leaf_88_core_clock),
    .D(_0222_),
    .Q(\dmmu0.page_table[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6962_ (.CLK(clknet_leaf_88_core_clock),
    .D(_0223_),
    .Q(\dmmu0.page_table[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6963_ (.CLK(clknet_leaf_88_core_clock),
    .D(_0224_),
    .Q(\dmmu0.page_table[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6964_ (.CLK(clknet_leaf_90_core_clock),
    .D(_0225_),
    .Q(\dmmu0.page_table[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6965_ (.CLK(clknet_leaf_87_core_clock),
    .D(_0226_),
    .Q(\dmmu0.page_table[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6966_ (.CLK(clknet_leaf_86_core_clock),
    .D(_0227_),
    .Q(\dmmu0.page_table[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6967_ (.CLK(clknet_leaf_89_core_clock),
    .D(_0228_),
    .Q(\dmmu0.page_table[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6968_ (.CLK(clknet_leaf_90_core_clock),
    .D(_0229_),
    .Q(\dmmu0.page_table[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6969_ (.CLK(clknet_leaf_86_core_clock),
    .D(_0230_),
    .Q(\dmmu0.page_table[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6970_ (.CLK(clknet_leaf_90_core_clock),
    .D(_0231_),
    .Q(\dmmu0.page_table[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6971_ (.CLK(clknet_leaf_90_core_clock),
    .D(_0232_),
    .Q(\dmmu0.page_table[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6972_ (.CLK(clknet_leaf_88_core_clock),
    .D(_0233_),
    .Q(\dmmu0.page_table[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6973_ (.CLK(clknet_leaf_0_core_clock),
    .D(_0234_),
    .Q(\dmmu0.page_table[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6974_ (.CLK(clknet_leaf_0_core_clock),
    .D(_0235_),
    .Q(\dmmu0.page_table[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6975_ (.CLK(clknet_leaf_0_core_clock),
    .D(_0236_),
    .Q(\dmmu0.page_table[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6976_ (.CLK(clknet_leaf_78_core_clock),
    .D(_0237_),
    .Q(\immu_0.high_addr_off[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6977_ (.CLK(clknet_leaf_11_core_clock),
    .D(_0238_),
    .Q(\immu_0.high_addr_off[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6978_ (.CLK(clknet_leaf_77_core_clock),
    .D(_0239_),
    .Q(\immu_0.high_addr_off[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6979_ (.CLK(clknet_leaf_57_core_clock),
    .D(_0240_),
    .Q(\immu_0.high_addr_off[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6980_ (.CLK(clknet_leaf_78_core_clock),
    .D(_0241_),
    .Q(\immu_0.high_addr_off[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6981_ (.CLK(clknet_leaf_78_core_clock),
    .D(_0242_),
    .Q(\immu_0.high_addr_off[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6982_ (.CLK(clknet_leaf_78_core_clock),
    .D(_0243_),
    .Q(\immu_0.high_addr_off[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6983_ (.CLK(clknet_leaf_78_core_clock),
    .D(_0244_),
    .Q(\immu_0.high_addr_off[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6984_ (.CLK(clknet_leaf_7_core_clock),
    .D(_0245_),
    .Q(\dmmu0.page_table[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6985_ (.CLK(clknet_leaf_7_core_clock),
    .D(_0246_),
    .Q(\dmmu0.page_table[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6986_ (.CLK(clknet_leaf_7_core_clock),
    .D(_0247_),
    .Q(\dmmu0.page_table[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6987_ (.CLK(clknet_leaf_7_core_clock),
    .D(_0248_),
    .Q(\dmmu0.page_table[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6988_ (.CLK(clknet_leaf_8_core_clock),
    .D(_0249_),
    .Q(\dmmu0.page_table[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6989_ (.CLK(clknet_leaf_7_core_clock),
    .D(_0250_),
    .Q(\dmmu0.page_table[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6990_ (.CLK(clknet_leaf_8_core_clock),
    .D(_0251_),
    .Q(\dmmu0.page_table[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6991_ (.CLK(clknet_leaf_9_core_clock),
    .D(_0252_),
    .Q(\dmmu0.page_table[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6992_ (.CLK(clknet_leaf_9_core_clock),
    .D(_0253_),
    .Q(\dmmu0.page_table[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6993_ (.CLK(clknet_leaf_5_core_clock),
    .D(_0254_),
    .Q(\dmmu0.page_table[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6994_ (.CLK(clknet_leaf_4_core_clock),
    .D(_0255_),
    .Q(\dmmu0.page_table[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6995_ (.CLK(clknet_leaf_1_core_clock),
    .D(_0256_),
    .Q(\dmmu0.page_table[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6996_ (.CLK(clknet_leaf_6_core_clock),
    .D(_0257_),
    .Q(\dmmu0.page_table[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6997_ (.CLK(clknet_leaf_62_core_clock),
    .D(_0258_),
    .Q(\icache_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__dfxtp_1 _6998_ (.CLK(clknet_leaf_39_core_clock),
    .D(_0259_),
    .Q(\immu_1.high_addr_off[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6999_ (.CLK(clknet_leaf_38_core_clock),
    .D(_0260_),
    .Q(\immu_1.high_addr_off[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7000_ (.CLK(clknet_leaf_37_core_clock),
    .D(_0261_),
    .Q(\immu_1.high_addr_off[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7001_ (.CLK(clknet_leaf_37_core_clock),
    .D(_0262_),
    .Q(\immu_1.high_addr_off[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7002_ (.CLK(clknet_leaf_37_core_clock),
    .D(_0263_),
    .Q(\immu_1.high_addr_off[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7003_ (.CLK(clknet_leaf_36_core_clock),
    .D(_0264_),
    .Q(\immu_1.high_addr_off[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7004_ (.CLK(clknet_leaf_36_core_clock),
    .D(_0265_),
    .Q(\immu_1.high_addr_off[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7005_ (.CLK(clknet_leaf_36_core_clock),
    .D(_0266_),
    .Q(\immu_1.high_addr_off[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7006_ (.CLK(clknet_leaf_80_core_clock),
    .D(_0267_),
    .Q(\dmmu0.page_table[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7007_ (.CLK(clknet_leaf_79_core_clock),
    .D(_0268_),
    .Q(\dmmu0.page_table[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7008_ (.CLK(clknet_leaf_79_core_clock),
    .D(_0269_),
    .Q(\dmmu0.page_table[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7009_ (.CLK(clknet_leaf_78_core_clock),
    .D(_0270_),
    .Q(\dmmu0.page_table[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7010_ (.CLK(clknet_leaf_78_core_clock),
    .D(_0271_),
    .Q(\dmmu0.page_table[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7011_ (.CLK(clknet_leaf_78_core_clock),
    .D(_0272_),
    .Q(\dmmu0.page_table[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7012_ (.CLK(clknet_leaf_78_core_clock),
    .D(_0273_),
    .Q(\dmmu0.page_table[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7013_ (.CLK(clknet_leaf_37_core_clock),
    .D(_0274_),
    .Q(\dmmu0.page_table[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7014_ (.CLK(clknet_leaf_38_core_clock),
    .D(_0275_),
    .Q(\dmmu0.page_table[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7015_ (.CLK(clknet_leaf_11_core_clock),
    .D(_0276_),
    .Q(\dmmu0.page_table[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7016_ (.CLK(clknet_leaf_17_core_clock),
    .D(_0277_),
    .Q(\dmmu0.page_table[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7017_ (.CLK(clknet_leaf_17_core_clock),
    .D(_0278_),
    .Q(\dmmu0.page_table[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7018_ (.CLK(clknet_leaf_4_core_clock),
    .D(_0279_),
    .Q(\dmmu0.page_table[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7019_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0280_),
    .Q(\dmmu0.page_table[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7020_ (.CLK(clknet_leaf_84_core_clock),
    .D(_0281_),
    .Q(\dmmu0.page_table[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7021_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0282_),
    .Q(\dmmu0.page_table[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7022_ (.CLK(clknet_leaf_83_core_clock),
    .D(_0283_),
    .Q(\dmmu0.page_table[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7023_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0284_),
    .Q(\dmmu0.page_table[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7024_ (.CLK(clknet_leaf_83_core_clock),
    .D(_0285_),
    .Q(\dmmu0.page_table[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7025_ (.CLK(clknet_leaf_83_core_clock),
    .D(_0286_),
    .Q(\dmmu0.page_table[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7026_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0287_),
    .Q(\dmmu0.page_table[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7027_ (.CLK(clknet_leaf_84_core_clock),
    .D(_0288_),
    .Q(\dmmu0.page_table[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7028_ (.CLK(clknet_leaf_82_core_clock),
    .D(_0289_),
    .Q(\dmmu0.page_table[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7029_ (.CLK(clknet_leaf_7_core_clock),
    .D(_0290_),
    .Q(\dmmu0.page_table[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7030_ (.CLK(clknet_leaf_7_core_clock),
    .D(_0291_),
    .Q(\dmmu0.page_table[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7031_ (.CLK(clknet_leaf_6_core_clock),
    .D(_0292_),
    .Q(\dmmu0.page_table[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7032_ (.CLK(clknet_leaf_13_core_clock),
    .D(_0293_),
    .Q(\dmmu0.page_table[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7033_ (.CLK(clknet_leaf_13_core_clock),
    .D(_0294_),
    .Q(\dmmu0.page_table[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7034_ (.CLK(clknet_leaf_13_core_clock),
    .D(_0295_),
    .Q(\dmmu0.page_table[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7035_ (.CLK(clknet_leaf_12_core_clock),
    .D(_0296_),
    .Q(\dmmu0.page_table[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7036_ (.CLK(clknet_leaf_11_core_clock),
    .D(_0297_),
    .Q(\dmmu0.page_table[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7037_ (.CLK(clknet_leaf_12_core_clock),
    .D(_0298_),
    .Q(\dmmu0.page_table[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7038_ (.CLK(clknet_leaf_9_core_clock),
    .D(_0299_),
    .Q(\dmmu0.page_table[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7039_ (.CLK(clknet_leaf_13_core_clock),
    .D(_0300_),
    .Q(\dmmu0.page_table[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7040_ (.CLK(clknet_leaf_12_core_clock),
    .D(_0301_),
    .Q(\dmmu0.page_table[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7041_ (.CLK(clknet_leaf_17_core_clock),
    .D(_0302_),
    .Q(\dmmu0.page_table[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7042_ (.CLK(clknet_leaf_17_core_clock),
    .D(_0303_),
    .Q(\dmmu0.page_table[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7043_ (.CLK(clknet_leaf_17_core_clock),
    .D(_0304_),
    .Q(\dmmu0.page_table[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7044_ (.CLK(clknet_leaf_4_core_clock),
    .D(_0305_),
    .Q(\dmmu0.page_table[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7045_ (.CLK(clknet_leaf_36_core_clock),
    .D(_0306_),
    .Q(\dmmu1.page_table[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7046_ (.CLK(clknet_leaf_32_core_clock),
    .D(_0307_),
    .Q(\dmmu1.page_table[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7047_ (.CLK(clknet_leaf_37_core_clock),
    .D(_0308_),
    .Q(\dmmu1.page_table[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7048_ (.CLK(clknet_leaf_37_core_clock),
    .D(_0309_),
    .Q(\dmmu1.page_table[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7049_ (.CLK(clknet_leaf_32_core_clock),
    .D(_0310_),
    .Q(\dmmu1.page_table[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7050_ (.CLK(clknet_leaf_36_core_clock),
    .D(_0311_),
    .Q(\dmmu1.page_table[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7051_ (.CLK(clknet_leaf_36_core_clock),
    .D(_0312_),
    .Q(\dmmu1.page_table[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7052_ (.CLK(clknet_leaf_32_core_clock),
    .D(_0313_),
    .Q(\dmmu1.page_table[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7053_ (.CLK(clknet_leaf_32_core_clock),
    .D(_0314_),
    .Q(\dmmu1.page_table[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7054_ (.CLK(clknet_leaf_31_core_clock),
    .D(_0315_),
    .Q(\dmmu1.page_table[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7055_ (.CLK(clknet_leaf_30_core_clock),
    .D(_0316_),
    .Q(\dmmu1.page_table[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7056_ (.CLK(clknet_leaf_31_core_clock),
    .D(_0317_),
    .Q(\dmmu1.page_table[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7057_ (.CLK(clknet_leaf_31_core_clock),
    .D(_0318_),
    .Q(\dmmu1.page_table[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7058_ (.CLK(clknet_leaf_80_core_clock),
    .D(_0319_),
    .Q(\dmmu0.page_table[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7059_ (.CLK(clknet_leaf_80_core_clock),
    .D(_0320_),
    .Q(\dmmu0.page_table[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7060_ (.CLK(clknet_leaf_79_core_clock),
    .D(_0321_),
    .Q(\dmmu0.page_table[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7061_ (.CLK(clknet_leaf_80_core_clock),
    .D(_0322_),
    .Q(\dmmu0.page_table[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7062_ (.CLK(clknet_leaf_10_core_clock),
    .D(_0323_),
    .Q(\dmmu0.page_table[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7063_ (.CLK(clknet_leaf_10_core_clock),
    .D(_0324_),
    .Q(\dmmu0.page_table[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7064_ (.CLK(clknet_leaf_10_core_clock),
    .D(_0325_),
    .Q(\dmmu0.page_table[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7065_ (.CLK(clknet_leaf_11_core_clock),
    .D(_0326_),
    .Q(\dmmu0.page_table[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7066_ (.CLK(clknet_leaf_10_core_clock),
    .D(_0327_),
    .Q(\dmmu0.page_table[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7067_ (.CLK(clknet_leaf_5_core_clock),
    .D(_0328_),
    .Q(\dmmu0.page_table[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7068_ (.CLK(clknet_leaf_4_core_clock),
    .D(_0329_),
    .Q(\dmmu0.page_table[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7069_ (.CLK(clknet_leaf_4_core_clock),
    .D(_0330_),
    .Q(\dmmu0.page_table[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7070_ (.CLK(clknet_leaf_4_core_clock),
    .D(_0331_),
    .Q(\dmmu0.page_table[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7071_ (.CLK(clknet_leaf_79_core_clock),
    .D(_0332_),
    .Q(\dmmu0.page_table[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7072_ (.CLK(clknet_leaf_79_core_clock),
    .D(_0333_),
    .Q(\dmmu0.page_table[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7073_ (.CLK(clknet_leaf_79_core_clock),
    .D(_0334_),
    .Q(\dmmu0.page_table[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7074_ (.CLK(clknet_leaf_79_core_clock),
    .D(_0335_),
    .Q(\dmmu0.page_table[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7075_ (.CLK(clknet_leaf_10_core_clock),
    .D(_0336_),
    .Q(\dmmu0.page_table[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7076_ (.CLK(clknet_leaf_79_core_clock),
    .D(_0337_),
    .Q(\dmmu0.page_table[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7077_ (.CLK(clknet_leaf_78_core_clock),
    .D(_0338_),
    .Q(\dmmu0.page_table[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7078_ (.CLK(clknet_leaf_11_core_clock),
    .D(_0339_),
    .Q(\dmmu0.page_table[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7079_ (.CLK(clknet_leaf_11_core_clock),
    .D(_0340_),
    .Q(\dmmu0.page_table[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7080_ (.CLK(clknet_leaf_11_core_clock),
    .D(_0341_),
    .Q(\dmmu0.page_table[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7081_ (.CLK(clknet_leaf_9_core_clock),
    .D(_0342_),
    .Q(\dmmu0.page_table[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7082_ (.CLK(clknet_leaf_5_core_clock),
    .D(_0343_),
    .Q(\dmmu0.page_table[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7083_ (.CLK(clknet_leaf_5_core_clock),
    .D(_0344_),
    .Q(\dmmu0.page_table[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7084_ (.CLK(clknet_leaf_93_core_clock),
    .D(_0345_),
    .Q(\dmmu0.long_off_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7085_ (.CLK(clknet_leaf_93_core_clock),
    .D(_0346_),
    .Q(\dmmu0.long_off_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7086_ (.CLK(clknet_leaf_0_core_clock),
    .D(_0347_),
    .Q(\dmmu0.long_off_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7087_ (.CLK(clknet_leaf_93_core_clock),
    .D(_0348_),
    .Q(\dmmu0.long_off_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7088_ (.CLK(clknet_leaf_2_core_clock),
    .D(_0349_),
    .Q(\dmmu0.long_off_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7089_ (.CLK(clknet_leaf_2_core_clock),
    .D(_0350_),
    .Q(\dmmu0.long_off_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7090_ (.CLK(clknet_leaf_2_core_clock),
    .D(_0351_),
    .Q(\dmmu0.long_off_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7091_ (.CLK(clknet_leaf_2_core_clock),
    .D(_0352_),
    .Q(\dmmu0.long_off_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7092_ (.CLK(clknet_leaf_35_core_clock),
    .D(_0353_),
    .Q(\dmmu1.page_table[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7093_ (.CLK(clknet_leaf_32_core_clock),
    .D(_0354_),
    .Q(\dmmu1.page_table[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7094_ (.CLK(clknet_leaf_11_core_clock),
    .D(_0355_),
    .Q(\dmmu1.page_table[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7095_ (.CLK(clknet_leaf_37_core_clock),
    .D(_0356_),
    .Q(\dmmu1.page_table[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7096_ (.CLK(clknet_leaf_32_core_clock),
    .D(_0357_),
    .Q(\dmmu1.page_table[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7097_ (.CLK(clknet_leaf_36_core_clock),
    .D(_0358_),
    .Q(\dmmu1.page_table[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7098_ (.CLK(clknet_leaf_35_core_clock),
    .D(_0359_),
    .Q(\dmmu1.page_table[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7099_ (.CLK(clknet_leaf_32_core_clock),
    .D(_0360_),
    .Q(\dmmu1.page_table[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7100_ (.CLK(clknet_leaf_32_core_clock),
    .D(_0361_),
    .Q(\dmmu1.page_table[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7101_ (.CLK(clknet_leaf_31_core_clock),
    .D(_0362_),
    .Q(\dmmu1.page_table[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7102_ (.CLK(clknet_leaf_30_core_clock),
    .D(_0363_),
    .Q(\dmmu1.page_table[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7103_ (.CLK(clknet_leaf_30_core_clock),
    .D(_0364_),
    .Q(\dmmu1.page_table[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7104_ (.CLK(clknet_leaf_30_core_clock),
    .D(_0365_),
    .Q(\dmmu1.page_table[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7105_ (.CLK(clknet_leaf_35_core_clock),
    .D(_0366_),
    .Q(\dmmu1.page_table[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7106_ (.CLK(clknet_leaf_32_core_clock),
    .D(_0367_),
    .Q(\dmmu1.page_table[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7107_ (.CLK(clknet_leaf_36_core_clock),
    .D(_0368_),
    .Q(\dmmu1.page_table[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7108_ (.CLK(clknet_leaf_37_core_clock),
    .D(_0369_),
    .Q(\dmmu1.page_table[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7109_ (.CLK(clknet_leaf_32_core_clock),
    .D(_0370_),
    .Q(\dmmu1.page_table[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7110_ (.CLK(clknet_leaf_35_core_clock),
    .D(_0371_),
    .Q(\dmmu1.page_table[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7111_ (.CLK(clknet_leaf_35_core_clock),
    .D(_0372_),
    .Q(\dmmu1.page_table[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7112_ (.CLK(clknet_leaf_32_core_clock),
    .D(_0373_),
    .Q(\dmmu1.page_table[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7113_ (.CLK(clknet_leaf_33_core_clock),
    .D(_0374_),
    .Q(\dmmu1.page_table[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7114_ (.CLK(clknet_leaf_31_core_clock),
    .D(_0375_),
    .Q(\dmmu1.page_table[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7115_ (.CLK(clknet_leaf_30_core_clock),
    .D(_0376_),
    .Q(\dmmu1.page_table[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7116_ (.CLK(clknet_leaf_30_core_clock),
    .D(_0377_),
    .Q(\dmmu1.page_table[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7117_ (.CLK(clknet_leaf_30_core_clock),
    .D(_0378_),
    .Q(\dmmu1.page_table[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7118_ (.CLK(clknet_leaf_14_core_clock),
    .D(_0379_),
    .Q(\dmmu1.page_table[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7119_ (.CLK(clknet_leaf_28_core_clock),
    .D(_0380_),
    .Q(\dmmu1.page_table[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7120_ (.CLK(clknet_leaf_14_core_clock),
    .D(_0381_),
    .Q(\dmmu1.page_table[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7121_ (.CLK(clknet_leaf_13_core_clock),
    .D(_0382_),
    .Q(\dmmu1.page_table[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7122_ (.CLK(clknet_leaf_34_core_clock),
    .D(_0383_),
    .Q(\dmmu1.page_table[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7123_ (.CLK(clknet_leaf_13_core_clock),
    .D(_0384_),
    .Q(\dmmu1.page_table[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7124_ (.CLK(clknet_leaf_34_core_clock),
    .D(_0385_),
    .Q(\dmmu1.page_table[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7125_ (.CLK(clknet_leaf_28_core_clock),
    .D(_0386_),
    .Q(\dmmu1.page_table[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7126_ (.CLK(clknet_leaf_33_core_clock),
    .D(_0387_),
    .Q(\dmmu1.page_table[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7127_ (.CLK(clknet_leaf_28_core_clock),
    .D(_0388_),
    .Q(\dmmu1.page_table[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7128_ (.CLK(clknet_leaf_29_core_clock),
    .D(_0389_),
    .Q(\dmmu1.page_table[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7129_ (.CLK(clknet_leaf_29_core_clock),
    .D(_0390_),
    .Q(\dmmu1.page_table[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7130_ (.CLK(clknet_leaf_29_core_clock),
    .D(_0391_),
    .Q(\dmmu1.page_table[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7131_ (.CLK(clknet_leaf_14_core_clock),
    .D(_0392_),
    .Q(\dmmu1.page_table[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7132_ (.CLK(clknet_leaf_34_core_clock),
    .D(_0393_),
    .Q(\dmmu1.page_table[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7133_ (.CLK(clknet_leaf_14_core_clock),
    .D(_0394_),
    .Q(\dmmu1.page_table[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7134_ (.CLK(clknet_leaf_13_core_clock),
    .D(_0395_),
    .Q(\dmmu1.page_table[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7135_ (.CLK(clknet_leaf_34_core_clock),
    .D(_0396_),
    .Q(\dmmu1.page_table[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7136_ (.CLK(clknet_leaf_13_core_clock),
    .D(_0397_),
    .Q(\dmmu1.page_table[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7137_ (.CLK(clknet_leaf_34_core_clock),
    .D(_0398_),
    .Q(\dmmu1.page_table[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7138_ (.CLK(clknet_leaf_28_core_clock),
    .D(_0399_),
    .Q(\dmmu1.page_table[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7139_ (.CLK(clknet_leaf_33_core_clock),
    .D(_0400_),
    .Q(\dmmu1.page_table[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7140_ (.CLK(clknet_leaf_29_core_clock),
    .D(_0401_),
    .Q(\dmmu1.page_table[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7141_ (.CLK(clknet_leaf_27_core_clock),
    .D(_0402_),
    .Q(\dmmu1.page_table[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7142_ (.CLK(clknet_leaf_29_core_clock),
    .D(_0403_),
    .Q(\dmmu1.page_table[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7143_ (.CLK(clknet_leaf_29_core_clock),
    .D(_0404_),
    .Q(\dmmu1.page_table[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7144_ (.CLK(clknet_leaf_34_core_clock),
    .D(_0405_),
    .Q(\dmmu1.page_table[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7145_ (.CLK(clknet_leaf_33_core_clock),
    .D(_0406_),
    .Q(\dmmu1.page_table[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7146_ (.CLK(clknet_leaf_14_core_clock),
    .D(_0407_),
    .Q(\dmmu1.page_table[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7147_ (.CLK(clknet_leaf_35_core_clock),
    .D(_0408_),
    .Q(\dmmu1.page_table[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7148_ (.CLK(clknet_leaf_34_core_clock),
    .D(_0409_),
    .Q(\dmmu1.page_table[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7149_ (.CLK(clknet_leaf_14_core_clock),
    .D(_0410_),
    .Q(\dmmu1.page_table[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7150_ (.CLK(clknet_leaf_35_core_clock),
    .D(_0411_),
    .Q(\dmmu1.page_table[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7151_ (.CLK(clknet_leaf_33_core_clock),
    .D(_0412_),
    .Q(\dmmu1.page_table[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7152_ (.CLK(clknet_leaf_33_core_clock),
    .D(_0413_),
    .Q(\dmmu1.page_table[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7153_ (.CLK(clknet_leaf_30_core_clock),
    .D(_0414_),
    .Q(\dmmu1.page_table[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7154_ (.CLK(clknet_leaf_29_core_clock),
    .D(_0415_),
    .Q(\dmmu1.page_table[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7155_ (.CLK(clknet_leaf_30_core_clock),
    .D(_0416_),
    .Q(\dmmu1.page_table[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7156_ (.CLK(clknet_leaf_29_core_clock),
    .D(_0417_),
    .Q(\dmmu1.page_table[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7157_ (.CLK(clknet_leaf_13_core_clock),
    .D(_0418_),
    .Q(\dmmu0.page_table[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7158_ (.CLK(clknet_leaf_12_core_clock),
    .D(_0419_),
    .Q(\dmmu0.page_table[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7159_ (.CLK(clknet_leaf_12_core_clock),
    .D(_0420_),
    .Q(\dmmu0.page_table[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7160_ (.CLK(clknet_leaf_12_core_clock),
    .D(_0421_),
    .Q(\dmmu0.page_table[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7161_ (.CLK(clknet_leaf_9_core_clock),
    .D(_0422_),
    .Q(\dmmu0.page_table[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7162_ (.CLK(clknet_leaf_11_core_clock),
    .D(_0423_),
    .Q(\dmmu0.page_table[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7163_ (.CLK(clknet_leaf_9_core_clock),
    .D(_0424_),
    .Q(\dmmu0.page_table[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7164_ (.CLK(clknet_leaf_9_core_clock),
    .D(_0425_),
    .Q(\dmmu0.page_table[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7165_ (.CLK(clknet_leaf_10_core_clock),
    .D(_0426_),
    .Q(\dmmu0.page_table[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7166_ (.CLK(clknet_leaf_17_core_clock),
    .D(_0427_),
    .Q(\dmmu0.page_table[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7167_ (.CLK(clknet_leaf_4_core_clock),
    .D(_0428_),
    .Q(\dmmu0.page_table[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7168_ (.CLK(clknet_leaf_4_core_clock),
    .D(_0429_),
    .Q(\dmmu0.page_table[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7169_ (.CLK(clknet_leaf_3_core_clock),
    .D(_0430_),
    .Q(\dmmu0.page_table[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7170_ (.CLK(clknet_leaf_35_core_clock),
    .D(_0431_),
    .Q(\dmmu1.page_table[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7171_ (.CLK(clknet_leaf_33_core_clock),
    .D(_0432_),
    .Q(\dmmu1.page_table[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7172_ (.CLK(clknet_leaf_37_core_clock),
    .D(_0433_),
    .Q(\dmmu1.page_table[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7173_ (.CLK(clknet_leaf_12_core_clock),
    .D(_0434_),
    .Q(\dmmu1.page_table[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7174_ (.CLK(clknet_leaf_35_core_clock),
    .D(_0435_),
    .Q(\dmmu1.page_table[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7175_ (.CLK(clknet_leaf_11_core_clock),
    .D(_0436_),
    .Q(\dmmu1.page_table[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7176_ (.CLK(clknet_leaf_34_core_clock),
    .D(_0437_),
    .Q(\dmmu1.page_table[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7177_ (.CLK(clknet_leaf_33_core_clock),
    .D(_0438_),
    .Q(\dmmu1.page_table[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7178_ (.CLK(clknet_leaf_33_core_clock),
    .D(_0439_),
    .Q(\dmmu1.page_table[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7179_ (.CLK(clknet_leaf_33_core_clock),
    .D(_0440_),
    .Q(\dmmu1.page_table[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7180_ (.CLK(clknet_leaf_29_core_clock),
    .D(_0441_),
    .Q(\dmmu1.page_table[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7181_ (.CLK(clknet_leaf_29_core_clock),
    .D(_0442_),
    .Q(\dmmu1.page_table[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7182_ (.CLK(clknet_leaf_29_core_clock),
    .D(_0443_),
    .Q(\dmmu1.page_table[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7183_ (.CLK(clknet_leaf_15_core_clock),
    .D(_0444_),
    .Q(\dmmu1.page_table[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7184_ (.CLK(clknet_leaf_28_core_clock),
    .D(_0445_),
    .Q(\dmmu1.page_table[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7185_ (.CLK(clknet_leaf_13_core_clock),
    .D(_0446_),
    .Q(\dmmu1.page_table[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7186_ (.CLK(clknet_leaf_16_core_clock),
    .D(_0447_),
    .Q(\dmmu1.page_table[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7187_ (.CLK(clknet_leaf_28_core_clock),
    .D(_0448_),
    .Q(\dmmu1.page_table[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7188_ (.CLK(clknet_leaf_14_core_clock),
    .D(_0449_),
    .Q(\dmmu1.page_table[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7189_ (.CLK(clknet_leaf_14_core_clock),
    .D(_0450_),
    .Q(\dmmu1.page_table[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7190_ (.CLK(clknet_leaf_15_core_clock),
    .D(_0451_),
    .Q(\dmmu1.page_table[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7191_ (.CLK(clknet_leaf_28_core_clock),
    .D(_0452_),
    .Q(\dmmu1.page_table[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7192_ (.CLK(clknet_leaf_27_core_clock),
    .D(_0453_),
    .Q(\dmmu1.page_table[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7193_ (.CLK(clknet_leaf_29_core_clock),
    .D(_0454_),
    .Q(\dmmu1.page_table[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7194_ (.CLK(clknet_leaf_27_core_clock),
    .D(_0455_),
    .Q(\dmmu1.page_table[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7195_ (.CLK(clknet_leaf_27_core_clock),
    .D(_0456_),
    .Q(\dmmu1.page_table[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7196_ (.CLK(clknet_leaf_16_core_clock),
    .D(_0457_),
    .Q(\dmmu1.page_table[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7197_ (.CLK(clknet_leaf_28_core_clock),
    .D(_0458_),
    .Q(\dmmu1.page_table[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7198_ (.CLK(clknet_leaf_16_core_clock),
    .D(_0459_),
    .Q(\dmmu1.page_table[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7199_ (.CLK(clknet_leaf_17_core_clock),
    .D(_0460_),
    .Q(\dmmu1.page_table[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7200_ (.CLK(clknet_leaf_22_core_clock),
    .D(_0461_),
    .Q(\dmmu1.page_table[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7201_ (.CLK(clknet_leaf_15_core_clock),
    .D(_0462_),
    .Q(\dmmu1.page_table[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7202_ (.CLK(clknet_leaf_15_core_clock),
    .D(_0463_),
    .Q(\dmmu1.page_table[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7203_ (.CLK(clknet_leaf_22_core_clock),
    .D(_0464_),
    .Q(\dmmu1.page_table[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7204_ (.CLK(clknet_leaf_23_core_clock),
    .D(_0465_),
    .Q(\dmmu1.page_table[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7205_ (.CLK(clknet_leaf_28_core_clock),
    .D(_0466_),
    .Q(\dmmu1.page_table[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7206_ (.CLK(clknet_leaf_27_core_clock),
    .D(_0467_),
    .Q(\dmmu1.page_table[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7207_ (.CLK(clknet_leaf_27_core_clock),
    .D(_0468_),
    .Q(\dmmu1.page_table[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7208_ (.CLK(clknet_leaf_27_core_clock),
    .D(_0469_),
    .Q(\dmmu1.page_table[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7209_ (.CLK(clknet_leaf_15_core_clock),
    .D(_0470_),
    .Q(\dmmu1.page_table[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7210_ (.CLK(clknet_leaf_23_core_clock),
    .D(_0471_),
    .Q(\dmmu1.page_table[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7211_ (.CLK(clknet_leaf_16_core_clock),
    .D(_0472_),
    .Q(\dmmu1.page_table[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7212_ (.CLK(clknet_leaf_16_core_clock),
    .D(_0473_),
    .Q(\dmmu1.page_table[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7213_ (.CLK(clknet_leaf_23_core_clock),
    .D(_0474_),
    .Q(\dmmu1.page_table[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7214_ (.CLK(clknet_leaf_15_core_clock),
    .D(_0475_),
    .Q(\dmmu1.page_table[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7215_ (.CLK(clknet_leaf_14_core_clock),
    .D(_0476_),
    .Q(\dmmu1.page_table[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7216_ (.CLK(clknet_leaf_22_core_clock),
    .D(_0477_),
    .Q(\dmmu1.page_table[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7217_ (.CLK(clknet_leaf_28_core_clock),
    .D(_0478_),
    .Q(\dmmu1.page_table[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7218_ (.CLK(clknet_leaf_28_core_clock),
    .D(_0479_),
    .Q(\dmmu1.page_table[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7219_ (.CLK(clknet_leaf_27_core_clock),
    .D(_0480_),
    .Q(\dmmu1.page_table[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7220_ (.CLK(clknet_leaf_27_core_clock),
    .D(_0481_),
    .Q(\dmmu1.page_table[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7221_ (.CLK(clknet_leaf_27_core_clock),
    .D(_0482_),
    .Q(\dmmu1.page_table[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7222_ (.CLK(clknet_leaf_16_core_clock),
    .D(_0483_),
    .Q(\dmmu1.page_table[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7223_ (.CLK(clknet_leaf_23_core_clock),
    .D(_0484_),
    .Q(\dmmu1.page_table[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7224_ (.CLK(clknet_leaf_17_core_clock),
    .D(_0485_),
    .Q(\dmmu1.page_table[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7225_ (.CLK(clknet_leaf_17_core_clock),
    .D(_0486_),
    .Q(\dmmu1.page_table[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7226_ (.CLK(clknet_leaf_22_core_clock),
    .D(_0487_),
    .Q(\dmmu1.page_table[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7227_ (.CLK(clknet_leaf_22_core_clock),
    .D(_0488_),
    .Q(\dmmu1.page_table[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7228_ (.CLK(clknet_leaf_22_core_clock),
    .D(_0489_),
    .Q(\dmmu1.page_table[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7229_ (.CLK(clknet_leaf_22_core_clock),
    .D(_0490_),
    .Q(\dmmu1.page_table[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7230_ (.CLK(clknet_leaf_23_core_clock),
    .D(_0491_),
    .Q(\dmmu1.page_table[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7231_ (.CLK(clknet_leaf_23_core_clock),
    .D(_0492_),
    .Q(\dmmu1.page_table[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7232_ (.CLK(clknet_leaf_27_core_clock),
    .D(_0493_),
    .Q(\dmmu1.page_table[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7233_ (.CLK(clknet_leaf_26_core_clock),
    .D(_0494_),
    .Q(\dmmu1.page_table[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7234_ (.CLK(clknet_leaf_26_core_clock),
    .D(_0495_),
    .Q(\dmmu1.page_table[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7235_ (.CLK(clknet_leaf_21_core_clock),
    .D(_0496_),
    .Q(\dmmu1.page_table[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7236_ (.CLK(clknet_leaf_24_core_clock),
    .D(_0497_),
    .Q(\dmmu1.page_table[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7237_ (.CLK(clknet_leaf_21_core_clock),
    .D(_0498_),
    .Q(\dmmu1.page_table[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7238_ (.CLK(clknet_leaf_20_core_clock),
    .D(_0499_),
    .Q(\dmmu1.page_table[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7239_ (.CLK(clknet_leaf_24_core_clock),
    .D(_0500_),
    .Q(\dmmu1.page_table[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7240_ (.CLK(clknet_leaf_20_core_clock),
    .D(_0501_),
    .Q(\dmmu1.page_table[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7241_ (.CLK(clknet_leaf_24_core_clock),
    .D(_0502_),
    .Q(\dmmu1.page_table[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7242_ (.CLK(clknet_leaf_21_core_clock),
    .D(_0503_),
    .Q(\dmmu1.page_table[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7243_ (.CLK(clknet_leaf_23_core_clock),
    .D(_0504_),
    .Q(\dmmu1.page_table[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7244_ (.CLK(clknet_leaf_23_core_clock),
    .D(_0505_),
    .Q(\dmmu1.page_table[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7245_ (.CLK(clknet_leaf_26_core_clock),
    .D(_0506_),
    .Q(\dmmu1.page_table[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7246_ (.CLK(clknet_leaf_26_core_clock),
    .D(_0507_),
    .Q(\dmmu1.page_table[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7247_ (.CLK(clknet_leaf_26_core_clock),
    .D(_0508_),
    .Q(\dmmu1.page_table[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7248_ (.CLK(clknet_leaf_20_core_clock),
    .D(_0509_),
    .Q(\dmmu1.page_table[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7249_ (.CLK(clknet_leaf_24_core_clock),
    .D(_0510_),
    .Q(\dmmu1.page_table[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7250_ (.CLK(clknet_leaf_20_core_clock),
    .D(_0511_),
    .Q(\dmmu1.page_table[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7251_ (.CLK(clknet_leaf_19_core_clock),
    .D(_0512_),
    .Q(\dmmu1.page_table[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7252_ (.CLK(clknet_leaf_24_core_clock),
    .D(_0513_),
    .Q(\dmmu1.page_table[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7253_ (.CLK(clknet_leaf_20_core_clock),
    .D(_0514_),
    .Q(\dmmu1.page_table[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7254_ (.CLK(clknet_leaf_21_core_clock),
    .D(_0515_),
    .Q(\dmmu1.page_table[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7255_ (.CLK(clknet_leaf_21_core_clock),
    .D(_0516_),
    .Q(\dmmu1.page_table[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7256_ (.CLK(clknet_leaf_24_core_clock),
    .D(_0517_),
    .Q(\dmmu1.page_table[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7257_ (.CLK(clknet_leaf_25_core_clock),
    .D(_0518_),
    .Q(\dmmu1.page_table[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7258_ (.CLK(clknet_leaf_25_core_clock),
    .D(_0519_),
    .Q(\dmmu1.page_table[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7259_ (.CLK(clknet_leaf_25_core_clock),
    .D(_0520_),
    .Q(\dmmu1.page_table[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7260_ (.CLK(clknet_leaf_25_core_clock),
    .D(_0521_),
    .Q(\dmmu1.page_table[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7261_ (.CLK(clknet_leaf_20_core_clock),
    .D(_0522_),
    .Q(\dmmu1.page_table[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7262_ (.CLK(clknet_leaf_25_core_clock),
    .D(_0523_),
    .Q(\dmmu1.page_table[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7263_ (.CLK(clknet_leaf_20_core_clock),
    .D(_0524_),
    .Q(\dmmu1.page_table[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7264_ (.CLK(clknet_leaf_19_core_clock),
    .D(_0525_),
    .Q(\dmmu1.page_table[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7265_ (.CLK(clknet_leaf_24_core_clock),
    .D(_0526_),
    .Q(\dmmu1.page_table[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7266_ (.CLK(clknet_leaf_20_core_clock),
    .D(_0527_),
    .Q(\dmmu1.page_table[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7267_ (.CLK(clknet_leaf_21_core_clock),
    .D(_0528_),
    .Q(\dmmu1.page_table[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7268_ (.CLK(clknet_leaf_21_core_clock),
    .D(_0529_),
    .Q(\dmmu1.page_table[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7269_ (.CLK(clknet_leaf_24_core_clock),
    .D(_0530_),
    .Q(\dmmu1.page_table[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7270_ (.CLK(clknet_leaf_25_core_clock),
    .D(_0531_),
    .Q(\dmmu1.page_table[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7271_ (.CLK(clknet_leaf_25_core_clock),
    .D(_0532_),
    .Q(\dmmu1.page_table[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7272_ (.CLK(clknet_leaf_26_core_clock),
    .D(_0533_),
    .Q(\dmmu1.page_table[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7273_ (.CLK(clknet_leaf_26_core_clock),
    .D(_0534_),
    .Q(\dmmu1.page_table[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7274_ (.CLK(clknet_leaf_20_core_clock),
    .D(_0535_),
    .Q(\dmmu1.page_table[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7275_ (.CLK(clknet_leaf_23_core_clock),
    .D(_0536_),
    .Q(\dmmu1.page_table[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7276_ (.CLK(clknet_leaf_22_core_clock),
    .D(_0537_),
    .Q(\dmmu1.page_table[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7277_ (.CLK(clknet_leaf_18_core_clock),
    .D(_0538_),
    .Q(\dmmu1.page_table[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7278_ (.CLK(clknet_leaf_21_core_clock),
    .D(_0539_),
    .Q(\dmmu1.page_table[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7279_ (.CLK(clknet_leaf_21_core_clock),
    .D(_0540_),
    .Q(\dmmu1.page_table[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7280_ (.CLK(clknet_leaf_21_core_clock),
    .D(_0541_),
    .Q(\dmmu1.page_table[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7281_ (.CLK(clknet_leaf_21_core_clock),
    .D(_0542_),
    .Q(\dmmu1.page_table[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7282_ (.CLK(clknet_leaf_24_core_clock),
    .D(_0543_),
    .Q(\dmmu1.page_table[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7283_ (.CLK(clknet_leaf_25_core_clock),
    .D(_0544_),
    .Q(\dmmu1.page_table[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7284_ (.CLK(clknet_leaf_26_core_clock),
    .D(_0545_),
    .Q(\dmmu1.page_table[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7285_ (.CLK(clknet_leaf_26_core_clock),
    .D(_0546_),
    .Q(\dmmu1.page_table[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7286_ (.CLK(clknet_leaf_26_core_clock),
    .D(_0547_),
    .Q(\dmmu1.page_table[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7287_ (.CLK(clknet_leaf_93_core_clock),
    .D(_0548_),
    .Q(\mem_dcache_arb.select ));
 sky130_fd_sc_hd__dfxtp_1 _7288_ (.CLK(clknet_leaf_3_core_clock),
    .D(_0549_),
    .Q(\mem_dcache_arb.req1_pending ));
 sky130_fd_sc_hd__dfxtp_1 _7289_ (.CLK(clknet_leaf_93_core_clock),
    .D(_0550_),
    .Q(\mem_dcache_arb.req0_pending ));
 sky130_fd_sc_hd__dfxtp_1 _7290_ (.CLK(clknet_leaf_92_core_clock),
    .D(_0551_),
    .Q(\mem_dcache_arb.transfer_active ));
 sky130_fd_sc_hd__dfxtp_1 _7291_ (.CLK(clknet_leaf_44_core_clock),
    .D(_0552_),
    .Q(\immu_1.page_table[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7292_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0553_),
    .Q(\immu_1.page_table[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7293_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0554_),
    .Q(\immu_1.page_table[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7294_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0555_),
    .Q(\immu_1.page_table[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7295_ (.CLK(clknet_leaf_44_core_clock),
    .D(_0556_),
    .Q(\immu_1.page_table[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7296_ (.CLK(clknet_leaf_44_core_clock),
    .D(_0557_),
    .Q(\immu_1.page_table[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7297_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0558_),
    .Q(\immu_1.page_table[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7298_ (.CLK(clknet_leaf_43_core_clock),
    .D(_0559_),
    .Q(\immu_1.page_table[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7299_ (.CLK(clknet_leaf_44_core_clock),
    .D(_0560_),
    .Q(\immu_1.page_table[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7300_ (.CLK(clknet_leaf_44_core_clock),
    .D(_0561_),
    .Q(\immu_1.page_table[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7301_ (.CLK(clknet_leaf_44_core_clock),
    .D(_0562_),
    .Q(\immu_1.page_table[8][10] ));
 sky130_fd_sc_hd__dfxtp_4 _7302_ (.CLK(clknet_leaf_62_core_clock),
    .D(_0563_),
    .Q(\inner_wb_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__dfxtp_1 _7303_ (.CLK(clknet_leaf_3_core_clock),
    .D(_0564_),
    .Q(\dmmu1.long_off_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7304_ (.CLK(clknet_leaf_3_core_clock),
    .D(_0565_),
    .Q(\dmmu1.long_off_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7305_ (.CLK(clknet_leaf_3_core_clock),
    .D(_0566_),
    .Q(\dmmu1.long_off_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7306_ (.CLK(clknet_leaf_18_core_clock),
    .D(_0567_),
    .Q(\dmmu1.long_off_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7307_ (.CLK(clknet_leaf_19_core_clock),
    .D(_0568_),
    .Q(\dmmu1.long_off_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7308_ (.CLK(clknet_leaf_19_core_clock),
    .D(_0569_),
    .Q(\dmmu1.long_off_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7309_ (.CLK(clknet_leaf_19_core_clock),
    .D(_0570_),
    .Q(\dmmu1.long_off_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7310_ (.CLK(clknet_leaf_3_core_clock),
    .D(_0571_),
    .Q(\dmmu1.long_off_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7311_ (.CLK(clknet_leaf_2_core_clock),
    .D(_0572_),
    .Q(\icore_sregs.c1_disable ));
 sky130_fd_sc_hd__conb_1 interconnect_inner_712 (.LO(net712));
 sky130_fd_sc_hd__conb_1 interconnect_inner_713 (.LO(net713));
 sky130_fd_sc_hd__conb_1 interconnect_inner_714 (.LO(net714));
 sky130_fd_sc_hd__conb_1 interconnect_inner_715 (.LO(net715));
 sky130_fd_sc_hd__conb_1 interconnect_inner_716 (.LO(net716));
 sky130_fd_sc_hd__conb_1 interconnect_inner_717 (.LO(net717));
 sky130_fd_sc_hd__conb_1 interconnect_inner_718 (.LO(net718));
 sky130_fd_sc_hd__conb_1 interconnect_inner_719 (.LO(net719));
 sky130_fd_sc_hd__conb_1 interconnect_inner_720 (.LO(net720));
 sky130_fd_sc_hd__conb_1 interconnect_inner_721 (.LO(net721));
 sky130_fd_sc_hd__conb_1 interconnect_inner_722 (.LO(net722));
 sky130_fd_sc_hd__conb_1 interconnect_inner_723 (.LO(net723));
 sky130_fd_sc_hd__conb_1 interconnect_inner_724 (.LO(net724));
 sky130_fd_sc_hd__conb_1 interconnect_inner_725 (.LO(net725));
 sky130_fd_sc_hd__conb_1 interconnect_inner_726 (.LO(net726));
 sky130_fd_sc_hd__conb_1 interconnect_inner_727 (.LO(net727));
 sky130_fd_sc_hd__conb_1 interconnect_inner_728 (.LO(net728));
 sky130_fd_sc_hd__conb_1 interconnect_inner_729 (.LO(net729));
 sky130_fd_sc_hd__conb_1 interconnect_inner_730 (.LO(net730));
 sky130_fd_sc_hd__conb_1 interconnect_inner_731 (.LO(net731));
 sky130_fd_sc_hd__conb_1 interconnect_inner_732 (.LO(net732));
 sky130_fd_sc_hd__conb_1 interconnect_inner_733 (.LO(net733));
 sky130_fd_sc_hd__conb_1 interconnect_inner_734 (.LO(net734));
 sky130_fd_sc_hd__conb_1 interconnect_inner_735 (.LO(net735));
 sky130_fd_sc_hd__conb_1 interconnect_inner_736 (.LO(net736));
 sky130_fd_sc_hd__conb_1 interconnect_inner_737 (.LO(net737));
 sky130_fd_sc_hd__conb_1 interconnect_inner_738 (.LO(net738));
 sky130_fd_sc_hd__conb_1 interconnect_inner_739 (.LO(net739));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_0_core_clock));
 sky130_fd_sc_hd__buf_2 _7341_ (.A(clknet_leaf_92_core_clock),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_1 _7342_ (.A(net384),
    .X(net406));
 sky130_fd_sc_hd__buf_4 _7343_ (.A(net386),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_1 _7344_ (.A(net407),
    .X(net410));
 sky130_fd_sc_hd__buf_2 _7345_ (.A(net277),
    .X(net429));
 sky130_fd_sc_hd__buf_2 _7346_ (.A(net288),
    .X(net440));
 sky130_fd_sc_hd__buf_2 _7347_ (.A(net299),
    .X(net451));
 sky130_fd_sc_hd__buf_2 _7348_ (.A(net302),
    .X(net454));
 sky130_fd_sc_hd__buf_2 _7349_ (.A(net303),
    .X(net455));
 sky130_fd_sc_hd__buf_2 _7350_ (.A(net304),
    .X(net456));
 sky130_fd_sc_hd__buf_2 _7351_ (.A(net305),
    .X(net457));
 sky130_fd_sc_hd__buf_2 _7352_ (.A(net306),
    .X(net458));
 sky130_fd_sc_hd__buf_2 _7353_ (.A(net307),
    .X(net459));
 sky130_fd_sc_hd__buf_2 _7354_ (.A(net308),
    .X(net460));
 sky130_fd_sc_hd__buf_2 _7355_ (.A(net278),
    .X(net430));
 sky130_fd_sc_hd__buf_2 _7356_ (.A(net279),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_2 _7357_ (.A(net280),
    .X(net432));
 sky130_fd_sc_hd__buf_2 _7358_ (.A(net281),
    .X(net433));
 sky130_fd_sc_hd__buf_2 _7359_ (.A(net282),
    .X(net434));
 sky130_fd_sc_hd__buf_2 _7360_ (.A(net283),
    .X(net435));
 sky130_fd_sc_hd__buf_2 _7361_ (.A(net284),
    .X(net436));
 sky130_fd_sc_hd__buf_2 _7362_ (.A(net285),
    .X(net437));
 sky130_fd_sc_hd__buf_2 _7363_ (.A(net286),
    .X(net438));
 sky130_fd_sc_hd__buf_2 _7364_ (.A(net287),
    .X(net439));
 sky130_fd_sc_hd__buf_2 _7365_ (.A(net289),
    .X(net441));
 sky130_fd_sc_hd__buf_2 _7366_ (.A(net290),
    .X(net442));
 sky130_fd_sc_hd__buf_2 _7367_ (.A(net291),
    .X(net443));
 sky130_fd_sc_hd__buf_2 _7368_ (.A(net292),
    .X(net444));
 sky130_fd_sc_hd__buf_2 _7369_ (.A(net293),
    .X(net445));
 sky130_fd_sc_hd__buf_2 _7370_ (.A(net294),
    .X(net446));
 sky130_fd_sc_hd__buf_2 _7371_ (.A(net295),
    .X(net447));
 sky130_fd_sc_hd__buf_2 _7372_ (.A(net296),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_2 _7373_ (.A(net297),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 _7374_ (.A(net298),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_2 _7375_ (.A(net300),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_2 _7376_ (.A(net301),
    .X(net453));
 sky130_fd_sc_hd__buf_2 _7377_ (.A(net276),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_1 _7378_ (.A(net710),
    .X(net462));
 sky130_fd_sc_hd__buf_2 _7379_ (.A(clknet_leaf_19_core_clock),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_1 _7380_ (.A(net407),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_1 _7381_ (.A(net408),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_1 _7382_ (.A(net408),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_2 _7383_ (.A(net331),
    .X(net486));
 sky130_fd_sc_hd__buf_2 _7384_ (.A(net342),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_1 _7385_ (.A(net353),
    .X(net508));
 sky130_fd_sc_hd__clkbuf_1 _7386_ (.A(net356),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_1 _7387_ (.A(net357),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_1 _7388_ (.A(net358),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_1 _7389_ (.A(net359),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_1 _7390_ (.A(net360),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_1 _7391_ (.A(net361),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_1 _7392_ (.A(net362),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_1 _7393_ (.A(net332),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_1 _7394_ (.A(net333),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_1 _7395_ (.A(net334),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_1 _7396_ (.A(net335),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_1 _7397_ (.A(net336),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_1 _7398_ (.A(net337),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_1 _7399_ (.A(net338),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_1 _7400_ (.A(net339),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_1 _7401_ (.A(net340),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_1 _7402_ (.A(net341),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_1 _7403_ (.A(net343),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_1 _7404_ (.A(net344),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_1 _7405_ (.A(net345),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_1 _7406_ (.A(net346),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_1 _7407_ (.A(net347),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_1 _7408_ (.A(net348),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_1 _7409_ (.A(net349),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_1 _7410_ (.A(net350),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_1 _7411_ (.A(net351),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_1 _7412_ (.A(net352),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_1 _7413_ (.A(net354),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_1 _7414_ (.A(net355),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_2 _7415_ (.A(net330),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_1 _7416_ (.A(net211),
    .X(net519));
 sky130_fd_sc_hd__buf_2 _7417_ (.A(clknet_leaf_92_core_clock),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_1 _7418_ (.A(net710),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_1 _7419_ (.A(net389),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_1 _7420_ (.A(net396),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_1 _7421_ (.A(net397),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_1 _7422_ (.A(net398),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_1 _7423_ (.A(net399),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_1 _7424_ (.A(net400),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_1 _7425_ (.A(net401),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_1 _7426_ (.A(net402),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_1 _7427_ (.A(net403),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_1 _7428_ (.A(net404),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_1 _7429_ (.A(net390),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_1 _7430_ (.A(net391),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_1 _7431_ (.A(net392),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_1 _7432_ (.A(net393),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_1 _7433_ (.A(net394),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_1 _7434_ (.A(net395),
    .X(net575));
 sky130_fd_sc_hd__buf_2 _7435_ (.A(clknet_opt_1_0_core_clock),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_1 _7436_ (.A(net59),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_1 _7437_ (.A(net66),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_1 _7438_ (.A(net67),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_1 _7439_ (.A(net68),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_1 _7440_ (.A(net69),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_1 _7441_ (.A(net70),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_1 _7442_ (.A(net71),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_1 _7443_ (.A(net72),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_1 _7444_ (.A(net73),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_1 _7445_ (.A(net74),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_1 _7446_ (.A(net60),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_1 _7447_ (.A(net61),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_1 _7448_ (.A(net62),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_1 _7449_ (.A(net63),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_1 _7450_ (.A(net64),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_1 _7451_ (.A(net65),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_1 _7452_ (.A(net4),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_1 _7453_ (.A(net75),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_1 _7454_ (.A(net58),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_1 _7455_ (.A(net710),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_1 _7456_ (.A(net389),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_1 _7457_ (.A(net396),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_1 _7458_ (.A(net397),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_1 _7459_ (.A(net398),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_1 _7460_ (.A(net399),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_1 _7461_ (.A(net400),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_1 _7462_ (.A(net401),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_1 _7463_ (.A(net402),
    .X(net621));
 sky130_fd_sc_hd__clkbuf_1 _7464_ (.A(net403),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_1 _7465_ (.A(net404),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_1 _7466_ (.A(net390),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_1 _7467_ (.A(net391),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_1 _7468_ (.A(net392),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_1 _7469_ (.A(net393),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_1 _7470_ (.A(net394),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_1 _7471_ (.A(net395),
    .X(net614));
 sky130_fd_sc_hd__buf_2 _7472_ (.A(clknet_opt_2_1_core_clock),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_1 _7473_ (.A(net164),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_1 _7474_ (.A(net171),
    .X(net632));
 sky130_fd_sc_hd__buf_2 _7475_ (.A(net172),
    .X(net633));
 sky130_fd_sc_hd__buf_2 _7476_ (.A(net173),
    .X(net634));
 sky130_fd_sc_hd__buf_2 _7477_ (.A(net174),
    .X(net635));
 sky130_fd_sc_hd__buf_2 _7478_ (.A(net175),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_2 _7479_ (.A(net176),
    .X(net637));
 sky130_fd_sc_hd__buf_2 _7480_ (.A(net177),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_2 _7481_ (.A(net178),
    .X(net639));
 sky130_fd_sc_hd__buf_2 _7482_ (.A(net179),
    .X(net640));
 sky130_fd_sc_hd__buf_2 _7483_ (.A(net165),
    .X(net626));
 sky130_fd_sc_hd__buf_2 _7484_ (.A(net166),
    .X(net627));
 sky130_fd_sc_hd__buf_2 _7485_ (.A(net167),
    .X(net628));
 sky130_fd_sc_hd__buf_2 _7486_ (.A(net168),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_2 _7487_ (.A(net169),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_2 _7488_ (.A(net170),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_1 _7489_ (.A(net109),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_1 _7490_ (.A(net180),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_1 _7491_ (.A(net163),
    .X(net643));
 sky130_fd_sc_hd__clkbuf_1 _7492_ (.A(net211),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_1 _7493_ (.A(net389),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_1 _7494_ (.A(net396),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_1 _7495_ (.A(net397),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_1 _7496_ (.A(net398),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_1 _7497_ (.A(net399),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_1 _7498_ (.A(net400),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_1 _7499_ (.A(net401),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_1 _7500_ (.A(net402),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_1 _7501_ (.A(net403),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_1 _7502_ (.A(net404),
    .X(net662));
 sky130_fd_sc_hd__clkbuf_1 _7503_ (.A(net390),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_1 _7504_ (.A(net391),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_1 _7505_ (.A(net392),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_1 _7506_ (.A(net393),
    .X(net651));
 sky130_fd_sc_hd__clkbuf_1 _7507_ (.A(net394),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_1 _7508_ (.A(net395),
    .X(net653));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(c0_o_c_data_page),
    .X(net1));
 sky130_fd_sc_hd__buf_6 input2 (.A(c0_o_c_instr_long),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(c0_o_c_instr_page),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(c0_o_icache_flush),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(c0_o_instr_long_addr[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(c0_o_instr_long_addr[1]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(c0_o_instr_long_addr[2]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(c0_o_instr_long_addr[3]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(c0_o_instr_long_addr[4]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input10 (.A(c0_o_instr_long_addr[5]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(c0_o_instr_long_addr[6]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(c0_o_instr_long_addr[7]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(c0_o_mem_addr[0]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(c0_o_mem_addr[10]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(c0_o_mem_addr[11]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(c0_o_mem_addr[12]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(c0_o_mem_addr[13]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(c0_o_mem_addr[14]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(c0_o_mem_addr[15]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(c0_o_mem_addr[1]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(c0_o_mem_addr[2]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(c0_o_mem_addr[3]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(c0_o_mem_addr[4]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(c0_o_mem_addr[5]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(c0_o_mem_addr[6]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(c0_o_mem_addr[7]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(c0_o_mem_addr[8]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(c0_o_mem_addr[9]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(c0_o_mem_data[0]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(c0_o_mem_data[10]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(c0_o_mem_data[11]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(c0_o_mem_data[12]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(c0_o_mem_data[13]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(c0_o_mem_data[14]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(c0_o_mem_data[15]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(c0_o_mem_data[1]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(c0_o_mem_data[2]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(c0_o_mem_data[3]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(c0_o_mem_data[4]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(c0_o_mem_data[5]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(c0_o_mem_data[6]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(c0_o_mem_data[7]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(c0_o_mem_data[8]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(c0_o_mem_data[9]),
    .X(net44));
 sky130_fd_sc_hd__dlymetal6s2s_1 input45 (.A(c0_o_mem_high_addr[0]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(c0_o_mem_high_addr[1]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(c0_o_mem_high_addr[2]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(c0_o_mem_high_addr[3]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(c0_o_mem_high_addr[4]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(c0_o_mem_high_addr[5]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(c0_o_mem_high_addr[6]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(c0_o_mem_high_addr[7]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(c0_o_mem_long_mode),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(c0_o_mem_req),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(c0_o_mem_sel[0]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(c0_o_mem_sel[1]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(c0_o_mem_we),
    .X(net57));
 sky130_fd_sc_hd__buf_2 input58 (.A(c0_o_req_active),
    .X(net58));
 sky130_fd_sc_hd__buf_2 input59 (.A(c0_o_req_addr[0]),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input60 (.A(c0_o_req_addr[10]),
    .X(net60));
 sky130_fd_sc_hd__buf_2 input61 (.A(c0_o_req_addr[11]),
    .X(net61));
 sky130_fd_sc_hd__buf_2 input62 (.A(c0_o_req_addr[12]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(c0_o_req_addr[13]),
    .X(net63));
 sky130_fd_sc_hd__buf_2 input64 (.A(c0_o_req_addr[14]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 input65 (.A(c0_o_req_addr[15]),
    .X(net65));
 sky130_fd_sc_hd__buf_2 input66 (.A(c0_o_req_addr[1]),
    .X(net66));
 sky130_fd_sc_hd__buf_2 input67 (.A(c0_o_req_addr[2]),
    .X(net67));
 sky130_fd_sc_hd__buf_2 input68 (.A(c0_o_req_addr[3]),
    .X(net68));
 sky130_fd_sc_hd__buf_2 input69 (.A(c0_o_req_addr[4]),
    .X(net69));
 sky130_fd_sc_hd__buf_2 input70 (.A(c0_o_req_addr[5]),
    .X(net70));
 sky130_fd_sc_hd__buf_2 input71 (.A(c0_o_req_addr[6]),
    .X(net71));
 sky130_fd_sc_hd__buf_2 input72 (.A(c0_o_req_addr[7]),
    .X(net72));
 sky130_fd_sc_hd__buf_2 input73 (.A(c0_o_req_addr[8]),
    .X(net73));
 sky130_fd_sc_hd__buf_2 input74 (.A(c0_o_req_addr[9]),
    .X(net74));
 sky130_fd_sc_hd__buf_2 input75 (.A(c0_o_req_ppl_submit),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 input76 (.A(c0_sr_bus_addr[0]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(c0_sr_bus_addr[10]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(c0_sr_bus_addr[11]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(c0_sr_bus_addr[12]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(c0_sr_bus_addr[13]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(c0_sr_bus_addr[14]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(c0_sr_bus_addr[15]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(c0_sr_bus_addr[1]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(c0_sr_bus_addr[2]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(c0_sr_bus_addr[3]),
    .X(net85));
 sky130_fd_sc_hd__dlymetal6s2s_1 input86 (.A(c0_sr_bus_addr[4]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(c0_sr_bus_addr[5]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(c0_sr_bus_addr[6]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(c0_sr_bus_addr[7]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(c0_sr_bus_addr[8]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(c0_sr_bus_addr[9]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(c0_sr_bus_data_o[0]),
    .X(net92));
 sky130_fd_sc_hd__buf_2 input93 (.A(c0_sr_bus_data_o[10]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 input94 (.A(c0_sr_bus_data_o[11]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 input95 (.A(c0_sr_bus_data_o[12]),
    .X(net95));
 sky130_fd_sc_hd__buf_6 input96 (.A(c0_sr_bus_data_o[1]),
    .X(net96));
 sky130_fd_sc_hd__buf_4 input97 (.A(c0_sr_bus_data_o[2]),
    .X(net97));
 sky130_fd_sc_hd__buf_4 input98 (.A(c0_sr_bus_data_o[3]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_4 input99 (.A(c0_sr_bus_data_o[4]),
    .X(net99));
 sky130_fd_sc_hd__buf_6 input100 (.A(c0_sr_bus_data_o[5]),
    .X(net100));
 sky130_fd_sc_hd__buf_4 input101 (.A(c0_sr_bus_data_o[6]),
    .X(net101));
 sky130_fd_sc_hd__buf_4 input102 (.A(c0_sr_bus_data_o[7]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 input103 (.A(c0_sr_bus_data_o[8]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 input104 (.A(c0_sr_bus_data_o[9]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(c0_sr_bus_we),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(c1_o_c_data_page),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 input107 (.A(c1_o_c_instr_long),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(c1_o_c_instr_page),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(c1_o_icache_flush),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(c1_o_instr_long_addr[0]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 input111 (.A(c1_o_instr_long_addr[1]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 input112 (.A(c1_o_instr_long_addr[2]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 input113 (.A(c1_o_instr_long_addr[3]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(c1_o_instr_long_addr[4]),
    .X(net114));
 sky130_fd_sc_hd__dlymetal6s2s_1 input115 (.A(c1_o_instr_long_addr[5]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(c1_o_instr_long_addr[6]),
    .X(net116));
 sky130_fd_sc_hd__dlymetal6s2s_1 input117 (.A(c1_o_instr_long_addr[7]),
    .X(net117));
 sky130_fd_sc_hd__buf_2 input118 (.A(c1_o_mem_addr[0]),
    .X(net118));
 sky130_fd_sc_hd__buf_2 input119 (.A(c1_o_mem_addr[10]),
    .X(net119));
 sky130_fd_sc_hd__buf_4 input120 (.A(c1_o_mem_addr[11]),
    .X(net120));
 sky130_fd_sc_hd__buf_4 input121 (.A(c1_o_mem_addr[12]),
    .X(net121));
 sky130_fd_sc_hd__buf_2 input122 (.A(c1_o_mem_addr[13]),
    .X(net122));
 sky130_fd_sc_hd__buf_4 input123 (.A(c1_o_mem_addr[14]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(c1_o_mem_addr[15]),
    .X(net124));
 sky130_fd_sc_hd__buf_2 input125 (.A(c1_o_mem_addr[1]),
    .X(net125));
 sky130_fd_sc_hd__buf_2 input126 (.A(c1_o_mem_addr[2]),
    .X(net126));
 sky130_fd_sc_hd__buf_2 input127 (.A(c1_o_mem_addr[3]),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(c1_o_mem_addr[4]),
    .X(net128));
 sky130_fd_sc_hd__buf_2 input129 (.A(c1_o_mem_addr[5]),
    .X(net129));
 sky130_fd_sc_hd__buf_2 input130 (.A(c1_o_mem_addr[6]),
    .X(net130));
 sky130_fd_sc_hd__buf_2 input131 (.A(c1_o_mem_addr[7]),
    .X(net131));
 sky130_fd_sc_hd__buf_2 input132 (.A(c1_o_mem_addr[8]),
    .X(net132));
 sky130_fd_sc_hd__buf_2 input133 (.A(c1_o_mem_addr[9]),
    .X(net133));
 sky130_fd_sc_hd__buf_2 input134 (.A(c1_o_mem_data[0]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(c1_o_mem_data[10]),
    .X(net135));
 sky130_fd_sc_hd__buf_2 input136 (.A(c1_o_mem_data[11]),
    .X(net136));
 sky130_fd_sc_hd__buf_2 input137 (.A(c1_o_mem_data[12]),
    .X(net137));
 sky130_fd_sc_hd__buf_2 input138 (.A(c1_o_mem_data[13]),
    .X(net138));
 sky130_fd_sc_hd__buf_2 input139 (.A(c1_o_mem_data[14]),
    .X(net139));
 sky130_fd_sc_hd__buf_2 input140 (.A(c1_o_mem_data[15]),
    .X(net140));
 sky130_fd_sc_hd__buf_2 input141 (.A(c1_o_mem_data[1]),
    .X(net141));
 sky130_fd_sc_hd__buf_2 input142 (.A(c1_o_mem_data[2]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(c1_o_mem_data[3]),
    .X(net143));
 sky130_fd_sc_hd__buf_2 input144 (.A(c1_o_mem_data[4]),
    .X(net144));
 sky130_fd_sc_hd__buf_2 input145 (.A(c1_o_mem_data[5]),
    .X(net145));
 sky130_fd_sc_hd__buf_2 input146 (.A(c1_o_mem_data[6]),
    .X(net146));
 sky130_fd_sc_hd__buf_2 input147 (.A(c1_o_mem_data[7]),
    .X(net147));
 sky130_fd_sc_hd__buf_2 input148 (.A(c1_o_mem_data[8]),
    .X(net148));
 sky130_fd_sc_hd__buf_2 input149 (.A(c1_o_mem_data[9]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 input150 (.A(c1_o_mem_high_addr[0]),
    .X(net150));
 sky130_fd_sc_hd__dlymetal6s2s_1 input151 (.A(c1_o_mem_high_addr[1]),
    .X(net151));
 sky130_fd_sc_hd__dlymetal6s2s_1 input152 (.A(c1_o_mem_high_addr[2]),
    .X(net152));
 sky130_fd_sc_hd__dlymetal6s2s_1 input153 (.A(c1_o_mem_high_addr[3]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(c1_o_mem_high_addr[4]),
    .X(net154));
 sky130_fd_sc_hd__dlymetal6s2s_1 input155 (.A(c1_o_mem_high_addr[5]),
    .X(net155));
 sky130_fd_sc_hd__dlymetal6s2s_1 input156 (.A(c1_o_mem_high_addr[6]),
    .X(net156));
 sky130_fd_sc_hd__dlymetal6s2s_1 input157 (.A(c1_o_mem_high_addr[7]),
    .X(net157));
 sky130_fd_sc_hd__buf_2 input158 (.A(c1_o_mem_long_mode),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(c1_o_mem_req),
    .X(net159));
 sky130_fd_sc_hd__buf_2 input160 (.A(c1_o_mem_sel[0]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 input161 (.A(c1_o_mem_sel[1]),
    .X(net161));
 sky130_fd_sc_hd__buf_2 input162 (.A(c1_o_mem_we),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 input163 (.A(c1_o_req_active),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 input164 (.A(c1_o_req_addr[0]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(c1_o_req_addr[10]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(c1_o_req_addr[11]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(c1_o_req_addr[12]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(c1_o_req_addr[13]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(c1_o_req_addr[14]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(c1_o_req_addr[15]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 input171 (.A(c1_o_req_addr[1]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 input172 (.A(c1_o_req_addr[2]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 input173 (.A(c1_o_req_addr[3]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(c1_o_req_addr[4]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(c1_o_req_addr[5]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(c1_o_req_addr[6]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(c1_o_req_addr[7]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(c1_o_req_addr[8]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(c1_o_req_addr[9]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input180 (.A(c1_o_req_ppl_submit),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 input181 (.A(c1_sr_bus_addr[0]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(c1_sr_bus_addr[10]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(c1_sr_bus_addr[11]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(c1_sr_bus_addr[12]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(c1_sr_bus_addr[13]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(c1_sr_bus_addr[14]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(c1_sr_bus_addr[15]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_4 input188 (.A(c1_sr_bus_addr[1]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_4 input189 (.A(c1_sr_bus_addr[2]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 input190 (.A(c1_sr_bus_addr[3]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(c1_sr_bus_addr[4]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(c1_sr_bus_addr[5]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(c1_sr_bus_addr[6]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(c1_sr_bus_addr[7]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(c1_sr_bus_addr[8]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(c1_sr_bus_addr[9]),
    .X(net196));
 sky130_fd_sc_hd__buf_4 input197 (.A(c1_sr_bus_data_o[0]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_4 input198 (.A(c1_sr_bus_data_o[10]),
    .X(net198));
 sky130_fd_sc_hd__buf_2 input199 (.A(c1_sr_bus_data_o[11]),
    .X(net199));
 sky130_fd_sc_hd__buf_2 input200 (.A(c1_sr_bus_data_o[12]),
    .X(net200));
 sky130_fd_sc_hd__buf_4 input201 (.A(c1_sr_bus_data_o[1]),
    .X(net201));
 sky130_fd_sc_hd__buf_2 input202 (.A(c1_sr_bus_data_o[2]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 input203 (.A(c1_sr_bus_data_o[3]),
    .X(net203));
 sky130_fd_sc_hd__buf_2 input204 (.A(c1_sr_bus_data_o[4]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_2 input205 (.A(c1_sr_bus_data_o[5]),
    .X(net205));
 sky130_fd_sc_hd__buf_2 input206 (.A(c1_sr_bus_data_o[6]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 input207 (.A(c1_sr_bus_data_o[7]),
    .X(net207));
 sky130_fd_sc_hd__buf_2 input208 (.A(c1_sr_bus_data_o[8]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_4 input209 (.A(c1_sr_bus_data_o[9]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 input210 (.A(c1_sr_bus_we),
    .X(net210));
 sky130_fd_sc_hd__buf_6 input211 (.A(core_reset),
    .X(net211));
 sky130_fd_sc_hd__buf_2 input212 (.A(dcache_mem_ack),
    .X(net212));
 sky130_fd_sc_hd__buf_2 input213 (.A(dcache_mem_exception),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 input214 (.A(dcache_mem_o_data[0]),
    .X(net214));
 sky130_fd_sc_hd__buf_4 input215 (.A(dcache_mem_o_data[10]),
    .X(net215));
 sky130_fd_sc_hd__buf_4 input216 (.A(dcache_mem_o_data[11]),
    .X(net216));
 sky130_fd_sc_hd__buf_4 input217 (.A(dcache_mem_o_data[12]),
    .X(net217));
 sky130_fd_sc_hd__buf_4 input218 (.A(dcache_mem_o_data[13]),
    .X(net218));
 sky130_fd_sc_hd__buf_4 input219 (.A(dcache_mem_o_data[14]),
    .X(net219));
 sky130_fd_sc_hd__buf_4 input220 (.A(dcache_mem_o_data[15]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 input221 (.A(dcache_mem_o_data[1]),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 input222 (.A(dcache_mem_o_data[2]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_4 input223 (.A(dcache_mem_o_data[3]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_4 input224 (.A(dcache_mem_o_data[4]),
    .X(net224));
 sky130_fd_sc_hd__buf_4 input225 (.A(dcache_mem_o_data[5]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 input226 (.A(dcache_mem_o_data[6]),
    .X(net226));
 sky130_fd_sc_hd__buf_4 input227 (.A(dcache_mem_o_data[7]),
    .X(net227));
 sky130_fd_sc_hd__buf_4 input228 (.A(dcache_mem_o_data[8]),
    .X(net228));
 sky130_fd_sc_hd__buf_4 input229 (.A(dcache_mem_o_data[9]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 input230 (.A(dcache_wb_4_burst),
    .X(net230));
 sky130_fd_sc_hd__buf_2 input231 (.A(dcache_wb_adr[0]),
    .X(net231));
 sky130_fd_sc_hd__buf_2 input232 (.A(dcache_wb_adr[10]),
    .X(net232));
 sky130_fd_sc_hd__buf_2 input233 (.A(dcache_wb_adr[11]),
    .X(net233));
 sky130_fd_sc_hd__buf_2 input234 (.A(dcache_wb_adr[12]),
    .X(net234));
 sky130_fd_sc_hd__buf_2 input235 (.A(dcache_wb_adr[13]),
    .X(net235));
 sky130_fd_sc_hd__buf_2 input236 (.A(dcache_wb_adr[14]),
    .X(net236));
 sky130_fd_sc_hd__buf_2 input237 (.A(dcache_wb_adr[15]),
    .X(net237));
 sky130_fd_sc_hd__buf_2 input238 (.A(dcache_wb_adr[16]),
    .X(net238));
 sky130_fd_sc_hd__buf_2 input239 (.A(dcache_wb_adr[17]),
    .X(net239));
 sky130_fd_sc_hd__buf_2 input240 (.A(dcache_wb_adr[18]),
    .X(net240));
 sky130_fd_sc_hd__buf_2 input241 (.A(dcache_wb_adr[19]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_4 input242 (.A(dcache_wb_adr[1]),
    .X(net242));
 sky130_fd_sc_hd__buf_2 input243 (.A(dcache_wb_adr[20]),
    .X(net243));
 sky130_fd_sc_hd__buf_2 input244 (.A(dcache_wb_adr[21]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_4 input245 (.A(dcache_wb_adr[22]),
    .X(net245));
 sky130_fd_sc_hd__buf_2 input246 (.A(dcache_wb_adr[23]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_4 input247 (.A(dcache_wb_adr[2]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_4 input248 (.A(dcache_wb_adr[3]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 input249 (.A(dcache_wb_adr[4]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_4 input250 (.A(dcache_wb_adr[5]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_4 input251 (.A(dcache_wb_adr[6]),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_4 input252 (.A(dcache_wb_adr[7]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_4 input253 (.A(dcache_wb_adr[8]),
    .X(net253));
 sky130_fd_sc_hd__buf_2 input254 (.A(dcache_wb_adr[9]),
    .X(net254));
 sky130_fd_sc_hd__buf_4 input255 (.A(dcache_wb_cyc),
    .X(net255));
 sky130_fd_sc_hd__buf_6 input256 (.A(dcache_wb_o_dat[0]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_1 input257 (.A(dcache_wb_o_dat[10]),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 input258 (.A(dcache_wb_o_dat[11]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 input259 (.A(dcache_wb_o_dat[12]),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 input260 (.A(dcache_wb_o_dat[13]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 input261 (.A(dcache_wb_o_dat[14]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 input262 (.A(dcache_wb_o_dat[15]),
    .X(net262));
 sky130_fd_sc_hd__buf_6 input263 (.A(dcache_wb_o_dat[1]),
    .X(net263));
 sky130_fd_sc_hd__buf_6 input264 (.A(dcache_wb_o_dat[2]),
    .X(net264));
 sky130_fd_sc_hd__buf_6 input265 (.A(dcache_wb_o_dat[3]),
    .X(net265));
 sky130_fd_sc_hd__buf_6 input266 (.A(dcache_wb_o_dat[4]),
    .X(net266));
 sky130_fd_sc_hd__buf_6 input267 (.A(dcache_wb_o_dat[5]),
    .X(net267));
 sky130_fd_sc_hd__buf_6 input268 (.A(dcache_wb_o_dat[6]),
    .X(net268));
 sky130_fd_sc_hd__buf_6 input269 (.A(dcache_wb_o_dat[7]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_8 input270 (.A(dcache_wb_o_dat[8]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 input271 (.A(dcache_wb_o_dat[9]),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_4 input272 (.A(dcache_wb_sel[0]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_4 input273 (.A(dcache_wb_sel[1]),
    .X(net273));
 sky130_fd_sc_hd__buf_2 input274 (.A(dcache_wb_stb),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 input275 (.A(dcache_wb_we),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_1 input276 (.A(ic0_mem_ack),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 input277 (.A(ic0_mem_data[0]),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 input278 (.A(ic0_mem_data[10]),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 input279 (.A(ic0_mem_data[11]),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 input280 (.A(ic0_mem_data[12]),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_1 input281 (.A(ic0_mem_data[13]),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 input282 (.A(ic0_mem_data[14]),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 input283 (.A(ic0_mem_data[15]),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 input284 (.A(ic0_mem_data[16]),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 input285 (.A(ic0_mem_data[17]),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 input286 (.A(ic0_mem_data[18]),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_1 input287 (.A(ic0_mem_data[19]),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 input288 (.A(ic0_mem_data[1]),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_1 input289 (.A(ic0_mem_data[20]),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 input290 (.A(ic0_mem_data[21]),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_1 input291 (.A(ic0_mem_data[22]),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_1 input292 (.A(ic0_mem_data[23]),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_1 input293 (.A(ic0_mem_data[24]),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_1 input294 (.A(ic0_mem_data[25]),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 input295 (.A(ic0_mem_data[26]),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_1 input296 (.A(ic0_mem_data[27]),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_1 input297 (.A(ic0_mem_data[28]),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_1 input298 (.A(ic0_mem_data[29]),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_1 input299 (.A(ic0_mem_data[2]),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 input300 (.A(ic0_mem_data[30]),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 input301 (.A(ic0_mem_data[31]),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_1 input302 (.A(ic0_mem_data[3]),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_1 input303 (.A(ic0_mem_data[4]),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 input304 (.A(ic0_mem_data[5]),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_1 input305 (.A(ic0_mem_data[6]),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 input306 (.A(ic0_mem_data[7]),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 input307 (.A(ic0_mem_data[8]),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_1 input308 (.A(ic0_mem_data[9]),
    .X(net308));
 sky130_fd_sc_hd__buf_2 input309 (.A(ic0_wb_adr[0]),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 input310 (.A(ic0_wb_adr[10]),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 input311 (.A(ic0_wb_adr[11]),
    .X(net311));
 sky130_fd_sc_hd__buf_6 input312 (.A(ic0_wb_adr[12]),
    .X(net312));
 sky130_fd_sc_hd__buf_4 input313 (.A(ic0_wb_adr[13]),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_2 input314 (.A(ic0_wb_adr[14]),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_4 input315 (.A(ic0_wb_adr[15]),
    .X(net315));
 sky130_fd_sc_hd__buf_2 input316 (.A(ic0_wb_adr[1]),
    .X(net316));
 sky130_fd_sc_hd__buf_2 input317 (.A(ic0_wb_adr[2]),
    .X(net317));
 sky130_fd_sc_hd__buf_2 input318 (.A(ic0_wb_adr[3]),
    .X(net318));
 sky130_fd_sc_hd__buf_2 input319 (.A(ic0_wb_adr[4]),
    .X(net319));
 sky130_fd_sc_hd__buf_2 input320 (.A(ic0_wb_adr[5]),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_2 input321 (.A(ic0_wb_adr[6]),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_2 input322 (.A(ic0_wb_adr[7]),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_2 input323 (.A(ic0_wb_adr[8]),
    .X(net323));
 sky130_fd_sc_hd__dlymetal6s2s_1 input324 (.A(ic0_wb_adr[9]),
    .X(net324));
 sky130_fd_sc_hd__buf_2 input325 (.A(ic0_wb_cyc),
    .X(net325));
 sky130_fd_sc_hd__buf_2 input326 (.A(ic0_wb_sel[0]),
    .X(net326));
 sky130_fd_sc_hd__buf_2 input327 (.A(ic0_wb_sel[1]),
    .X(net327));
 sky130_fd_sc_hd__buf_2 input328 (.A(ic0_wb_stb),
    .X(net328));
 sky130_fd_sc_hd__buf_2 input329 (.A(ic0_wb_we),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_1 input330 (.A(ic1_mem_ack),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 input331 (.A(ic1_mem_data[0]),
    .X(net331));
 sky130_fd_sc_hd__buf_2 input332 (.A(ic1_mem_data[10]),
    .X(net332));
 sky130_fd_sc_hd__buf_2 input333 (.A(ic1_mem_data[11]),
    .X(net333));
 sky130_fd_sc_hd__buf_2 input334 (.A(ic1_mem_data[12]),
    .X(net334));
 sky130_fd_sc_hd__buf_2 input335 (.A(ic1_mem_data[13]),
    .X(net335));
 sky130_fd_sc_hd__buf_2 input336 (.A(ic1_mem_data[14]),
    .X(net336));
 sky130_fd_sc_hd__buf_2 input337 (.A(ic1_mem_data[15]),
    .X(net337));
 sky130_fd_sc_hd__buf_2 input338 (.A(ic1_mem_data[16]),
    .X(net338));
 sky130_fd_sc_hd__buf_2 input339 (.A(ic1_mem_data[17]),
    .X(net339));
 sky130_fd_sc_hd__buf_2 input340 (.A(ic1_mem_data[18]),
    .X(net340));
 sky130_fd_sc_hd__buf_2 input341 (.A(ic1_mem_data[19]),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_1 input342 (.A(ic1_mem_data[1]),
    .X(net342));
 sky130_fd_sc_hd__buf_2 input343 (.A(ic1_mem_data[20]),
    .X(net343));
 sky130_fd_sc_hd__buf_2 input344 (.A(ic1_mem_data[21]),
    .X(net344));
 sky130_fd_sc_hd__buf_2 input345 (.A(ic1_mem_data[22]),
    .X(net345));
 sky130_fd_sc_hd__buf_2 input346 (.A(ic1_mem_data[23]),
    .X(net346));
 sky130_fd_sc_hd__buf_2 input347 (.A(ic1_mem_data[24]),
    .X(net347));
 sky130_fd_sc_hd__buf_2 input348 (.A(ic1_mem_data[25]),
    .X(net348));
 sky130_fd_sc_hd__buf_2 input349 (.A(ic1_mem_data[26]),
    .X(net349));
 sky130_fd_sc_hd__buf_2 input350 (.A(ic1_mem_data[27]),
    .X(net350));
 sky130_fd_sc_hd__buf_2 input351 (.A(ic1_mem_data[28]),
    .X(net351));
 sky130_fd_sc_hd__buf_2 input352 (.A(ic1_mem_data[29]),
    .X(net352));
 sky130_fd_sc_hd__buf_2 input353 (.A(ic1_mem_data[2]),
    .X(net353));
 sky130_fd_sc_hd__buf_2 input354 (.A(ic1_mem_data[30]),
    .X(net354));
 sky130_fd_sc_hd__buf_2 input355 (.A(ic1_mem_data[31]),
    .X(net355));
 sky130_fd_sc_hd__buf_2 input356 (.A(ic1_mem_data[3]),
    .X(net356));
 sky130_fd_sc_hd__buf_2 input357 (.A(ic1_mem_data[4]),
    .X(net357));
 sky130_fd_sc_hd__buf_2 input358 (.A(ic1_mem_data[5]),
    .X(net358));
 sky130_fd_sc_hd__buf_2 input359 (.A(ic1_mem_data[6]),
    .X(net359));
 sky130_fd_sc_hd__buf_2 input360 (.A(ic1_mem_data[7]),
    .X(net360));
 sky130_fd_sc_hd__buf_2 input361 (.A(ic1_mem_data[8]),
    .X(net361));
 sky130_fd_sc_hd__buf_2 input362 (.A(ic1_mem_data[9]),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_1 input363 (.A(ic1_wb_adr[0]),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 input364 (.A(ic1_wb_adr[10]),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 input365 (.A(ic1_wb_adr[11]),
    .X(net365));
 sky130_fd_sc_hd__buf_2 input366 (.A(ic1_wb_adr[12]),
    .X(net366));
 sky130_fd_sc_hd__buf_4 input367 (.A(ic1_wb_adr[13]),
    .X(net367));
 sky130_fd_sc_hd__buf_2 input368 (.A(ic1_wb_adr[14]),
    .X(net368));
 sky130_fd_sc_hd__buf_4 input369 (.A(ic1_wb_adr[15]),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 input370 (.A(ic1_wb_adr[1]),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_1 input371 (.A(ic1_wb_adr[2]),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 input372 (.A(ic1_wb_adr[3]),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_1 input373 (.A(ic1_wb_adr[4]),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_1 input374 (.A(ic1_wb_adr[5]),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_1 input375 (.A(ic1_wb_adr[6]),
    .X(net375));
 sky130_fd_sc_hd__dlymetal6s2s_1 input376 (.A(ic1_wb_adr[7]),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_2 input377 (.A(ic1_wb_adr[8]),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_2 input378 (.A(ic1_wb_adr[9]),
    .X(net378));
 sky130_fd_sc_hd__dlymetal6s2s_1 input379 (.A(ic1_wb_cyc),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_1 input380 (.A(ic1_wb_sel[0]),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_1 input381 (.A(ic1_wb_sel[1]),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 input382 (.A(ic1_wb_stb),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_1 input383 (.A(ic1_wb_we),
    .X(net383));
 sky130_fd_sc_hd__buf_4 input384 (.A(inner_disable),
    .X(net384));
 sky130_fd_sc_hd__buf_6 input385 (.A(inner_embed_mode),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_1 input386 (.A(inner_ext_irq),
    .X(net386));
 sky130_fd_sc_hd__buf_8 input387 (.A(inner_wb_ack),
    .X(net387));
 sky130_fd_sc_hd__buf_8 input388 (.A(inner_wb_err),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_16 input389 (.A(inner_wb_i_dat[0]),
    .X(net389));
 sky130_fd_sc_hd__buf_8 input390 (.A(inner_wb_i_dat[10]),
    .X(net390));
 sky130_fd_sc_hd__buf_6 input391 (.A(inner_wb_i_dat[11]),
    .X(net391));
 sky130_fd_sc_hd__buf_6 input392 (.A(inner_wb_i_dat[12]),
    .X(net392));
 sky130_fd_sc_hd__buf_6 input393 (.A(inner_wb_i_dat[13]),
    .X(net393));
 sky130_fd_sc_hd__buf_6 input394 (.A(inner_wb_i_dat[14]),
    .X(net394));
 sky130_fd_sc_hd__buf_6 input395 (.A(inner_wb_i_dat[15]),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_16 input396 (.A(inner_wb_i_dat[1]),
    .X(net396));
 sky130_fd_sc_hd__buf_8 input397 (.A(inner_wb_i_dat[2]),
    .X(net397));
 sky130_fd_sc_hd__buf_8 input398 (.A(inner_wb_i_dat[3]),
    .X(net398));
 sky130_fd_sc_hd__buf_8 input399 (.A(inner_wb_i_dat[4]),
    .X(net399));
 sky130_fd_sc_hd__buf_8 input400 (.A(inner_wb_i_dat[5]),
    .X(net400));
 sky130_fd_sc_hd__buf_8 input401 (.A(inner_wb_i_dat[6]),
    .X(net401));
 sky130_fd_sc_hd__buf_8 input402 (.A(inner_wb_i_dat[7]),
    .X(net402));
 sky130_fd_sc_hd__buf_8 input403 (.A(inner_wb_i_dat[8]),
    .X(net403));
 sky130_fd_sc_hd__buf_8 input404 (.A(inner_wb_i_dat[9]),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_1 output405 (.A(net405),
    .X(c0_clk));
 sky130_fd_sc_hd__buf_2 output406 (.A(net406),
    .X(c0_disable));
 sky130_fd_sc_hd__buf_2 output407 (.A(net407),
    .X(c0_i_core_int_sreg[0]));
 sky130_fd_sc_hd__buf_2 output408 (.A(net408),
    .X(c0_i_core_int_sreg[1]));
 sky130_fd_sc_hd__buf_2 output409 (.A(net409),
    .X(c0_i_irq));
 sky130_fd_sc_hd__buf_2 output410 (.A(net410),
    .X(c0_i_mc_core_int));
 sky130_fd_sc_hd__buf_2 output411 (.A(net411),
    .X(c0_i_mem_ack));
 sky130_fd_sc_hd__buf_2 output412 (.A(net412),
    .X(c0_i_mem_data[0]));
 sky130_fd_sc_hd__buf_2 output413 (.A(net413),
    .X(c0_i_mem_data[10]));
 sky130_fd_sc_hd__buf_2 output414 (.A(net414),
    .X(c0_i_mem_data[11]));
 sky130_fd_sc_hd__buf_2 output415 (.A(net415),
    .X(c0_i_mem_data[12]));
 sky130_fd_sc_hd__buf_2 output416 (.A(net416),
    .X(c0_i_mem_data[13]));
 sky130_fd_sc_hd__buf_2 output417 (.A(net417),
    .X(c0_i_mem_data[14]));
 sky130_fd_sc_hd__buf_2 output418 (.A(net418),
    .X(c0_i_mem_data[15]));
 sky130_fd_sc_hd__buf_2 output419 (.A(net419),
    .X(c0_i_mem_data[1]));
 sky130_fd_sc_hd__buf_2 output420 (.A(net420),
    .X(c0_i_mem_data[2]));
 sky130_fd_sc_hd__buf_2 output421 (.A(net421),
    .X(c0_i_mem_data[3]));
 sky130_fd_sc_hd__buf_2 output422 (.A(net422),
    .X(c0_i_mem_data[4]));
 sky130_fd_sc_hd__buf_2 output423 (.A(net423),
    .X(c0_i_mem_data[5]));
 sky130_fd_sc_hd__buf_2 output424 (.A(net424),
    .X(c0_i_mem_data[6]));
 sky130_fd_sc_hd__buf_2 output425 (.A(net425),
    .X(c0_i_mem_data[7]));
 sky130_fd_sc_hd__buf_2 output426 (.A(net426),
    .X(c0_i_mem_data[8]));
 sky130_fd_sc_hd__buf_2 output427 (.A(net427),
    .X(c0_i_mem_data[9]));
 sky130_fd_sc_hd__buf_2 output428 (.A(net428),
    .X(c0_i_mem_exception));
 sky130_fd_sc_hd__buf_2 output429 (.A(net429),
    .X(c0_i_req_data[0]));
 sky130_fd_sc_hd__buf_2 output430 (.A(net430),
    .X(c0_i_req_data[10]));
 sky130_fd_sc_hd__buf_2 output431 (.A(net431),
    .X(c0_i_req_data[11]));
 sky130_fd_sc_hd__buf_2 output432 (.A(net432),
    .X(c0_i_req_data[12]));
 sky130_fd_sc_hd__buf_2 output433 (.A(net433),
    .X(c0_i_req_data[13]));
 sky130_fd_sc_hd__buf_2 output434 (.A(net434),
    .X(c0_i_req_data[14]));
 sky130_fd_sc_hd__buf_2 output435 (.A(net435),
    .X(c0_i_req_data[15]));
 sky130_fd_sc_hd__buf_2 output436 (.A(net436),
    .X(c0_i_req_data[16]));
 sky130_fd_sc_hd__buf_2 output437 (.A(net437),
    .X(c0_i_req_data[17]));
 sky130_fd_sc_hd__buf_2 output438 (.A(net438),
    .X(c0_i_req_data[18]));
 sky130_fd_sc_hd__buf_2 output439 (.A(net439),
    .X(c0_i_req_data[19]));
 sky130_fd_sc_hd__buf_2 output440 (.A(net440),
    .X(c0_i_req_data[1]));
 sky130_fd_sc_hd__buf_2 output441 (.A(net441),
    .X(c0_i_req_data[20]));
 sky130_fd_sc_hd__buf_2 output442 (.A(net442),
    .X(c0_i_req_data[21]));
 sky130_fd_sc_hd__buf_2 output443 (.A(net443),
    .X(c0_i_req_data[22]));
 sky130_fd_sc_hd__buf_2 output444 (.A(net444),
    .X(c0_i_req_data[23]));
 sky130_fd_sc_hd__buf_2 output445 (.A(net445),
    .X(c0_i_req_data[24]));
 sky130_fd_sc_hd__buf_2 output446 (.A(net446),
    .X(c0_i_req_data[25]));
 sky130_fd_sc_hd__buf_2 output447 (.A(net447),
    .X(c0_i_req_data[26]));
 sky130_fd_sc_hd__buf_2 output448 (.A(net448),
    .X(c0_i_req_data[27]));
 sky130_fd_sc_hd__buf_2 output449 (.A(net449),
    .X(c0_i_req_data[28]));
 sky130_fd_sc_hd__buf_2 output450 (.A(net450),
    .X(c0_i_req_data[29]));
 sky130_fd_sc_hd__buf_2 output451 (.A(net451),
    .X(c0_i_req_data[2]));
 sky130_fd_sc_hd__buf_2 output452 (.A(net452),
    .X(c0_i_req_data[30]));
 sky130_fd_sc_hd__buf_2 output453 (.A(net453),
    .X(c0_i_req_data[31]));
 sky130_fd_sc_hd__buf_2 output454 (.A(net454),
    .X(c0_i_req_data[3]));
 sky130_fd_sc_hd__buf_2 output455 (.A(net455),
    .X(c0_i_req_data[4]));
 sky130_fd_sc_hd__buf_2 output456 (.A(net456),
    .X(c0_i_req_data[5]));
 sky130_fd_sc_hd__buf_2 output457 (.A(net457),
    .X(c0_i_req_data[6]));
 sky130_fd_sc_hd__buf_2 output458 (.A(net458),
    .X(c0_i_req_data[7]));
 sky130_fd_sc_hd__buf_2 output459 (.A(net459),
    .X(c0_i_req_data[8]));
 sky130_fd_sc_hd__buf_2 output460 (.A(net460),
    .X(c0_i_req_data[9]));
 sky130_fd_sc_hd__buf_2 output461 (.A(net461),
    .X(c0_i_req_data_valid));
 sky130_fd_sc_hd__buf_2 output462 (.A(net462),
    .X(c0_rst));
 sky130_fd_sc_hd__clkbuf_1 output463 (.A(net463),
    .X(c1_clk));
 sky130_fd_sc_hd__buf_2 output464 (.A(net464),
    .X(c1_disable));
 sky130_fd_sc_hd__buf_2 output465 (.A(net465),
    .X(c1_i_core_int_sreg[0]));
 sky130_fd_sc_hd__buf_2 output466 (.A(net466),
    .X(c1_i_core_int_sreg[1]));
 sky130_fd_sc_hd__buf_2 output467 (.A(net467),
    .X(c1_i_mc_core_int));
 sky130_fd_sc_hd__buf_2 output468 (.A(net468),
    .X(c1_i_mem_ack));
 sky130_fd_sc_hd__buf_2 output469 (.A(net469),
    .X(c1_i_mem_data[0]));
 sky130_fd_sc_hd__buf_2 output470 (.A(net470),
    .X(c1_i_mem_data[10]));
 sky130_fd_sc_hd__buf_2 output471 (.A(net471),
    .X(c1_i_mem_data[11]));
 sky130_fd_sc_hd__buf_2 output472 (.A(net472),
    .X(c1_i_mem_data[12]));
 sky130_fd_sc_hd__buf_2 output473 (.A(net473),
    .X(c1_i_mem_data[13]));
 sky130_fd_sc_hd__buf_2 output474 (.A(net474),
    .X(c1_i_mem_data[14]));
 sky130_fd_sc_hd__buf_2 output475 (.A(net475),
    .X(c1_i_mem_data[15]));
 sky130_fd_sc_hd__buf_2 output476 (.A(net476),
    .X(c1_i_mem_data[1]));
 sky130_fd_sc_hd__buf_2 output477 (.A(net477),
    .X(c1_i_mem_data[2]));
 sky130_fd_sc_hd__buf_2 output478 (.A(net478),
    .X(c1_i_mem_data[3]));
 sky130_fd_sc_hd__buf_2 output479 (.A(net479),
    .X(c1_i_mem_data[4]));
 sky130_fd_sc_hd__buf_2 output480 (.A(net480),
    .X(c1_i_mem_data[5]));
 sky130_fd_sc_hd__buf_2 output481 (.A(net481),
    .X(c1_i_mem_data[6]));
 sky130_fd_sc_hd__buf_2 output482 (.A(net482),
    .X(c1_i_mem_data[7]));
 sky130_fd_sc_hd__buf_2 output483 (.A(net483),
    .X(c1_i_mem_data[8]));
 sky130_fd_sc_hd__buf_2 output484 (.A(net484),
    .X(c1_i_mem_data[9]));
 sky130_fd_sc_hd__buf_2 output485 (.A(net485),
    .X(c1_i_mem_exception));
 sky130_fd_sc_hd__buf_2 output486 (.A(net486),
    .X(c1_i_req_data[0]));
 sky130_fd_sc_hd__buf_2 output487 (.A(net487),
    .X(c1_i_req_data[10]));
 sky130_fd_sc_hd__buf_2 output488 (.A(net488),
    .X(c1_i_req_data[11]));
 sky130_fd_sc_hd__buf_2 output489 (.A(net489),
    .X(c1_i_req_data[12]));
 sky130_fd_sc_hd__buf_2 output490 (.A(net490),
    .X(c1_i_req_data[13]));
 sky130_fd_sc_hd__buf_2 output491 (.A(net491),
    .X(c1_i_req_data[14]));
 sky130_fd_sc_hd__buf_2 output492 (.A(net492),
    .X(c1_i_req_data[15]));
 sky130_fd_sc_hd__buf_2 output493 (.A(net493),
    .X(c1_i_req_data[16]));
 sky130_fd_sc_hd__buf_2 output494 (.A(net494),
    .X(c1_i_req_data[17]));
 sky130_fd_sc_hd__buf_2 output495 (.A(net495),
    .X(c1_i_req_data[18]));
 sky130_fd_sc_hd__buf_2 output496 (.A(net496),
    .X(c1_i_req_data[19]));
 sky130_fd_sc_hd__buf_2 output497 (.A(net497),
    .X(c1_i_req_data[1]));
 sky130_fd_sc_hd__buf_2 output498 (.A(net498),
    .X(c1_i_req_data[20]));
 sky130_fd_sc_hd__buf_2 output499 (.A(net499),
    .X(c1_i_req_data[21]));
 sky130_fd_sc_hd__buf_2 output500 (.A(net500),
    .X(c1_i_req_data[22]));
 sky130_fd_sc_hd__buf_2 output501 (.A(net501),
    .X(c1_i_req_data[23]));
 sky130_fd_sc_hd__buf_2 output502 (.A(net502),
    .X(c1_i_req_data[24]));
 sky130_fd_sc_hd__buf_2 output503 (.A(net503),
    .X(c1_i_req_data[25]));
 sky130_fd_sc_hd__buf_2 output504 (.A(net504),
    .X(c1_i_req_data[26]));
 sky130_fd_sc_hd__buf_2 output505 (.A(net505),
    .X(c1_i_req_data[27]));
 sky130_fd_sc_hd__buf_2 output506 (.A(net506),
    .X(c1_i_req_data[28]));
 sky130_fd_sc_hd__buf_2 output507 (.A(net507),
    .X(c1_i_req_data[29]));
 sky130_fd_sc_hd__buf_2 output508 (.A(net508),
    .X(c1_i_req_data[2]));
 sky130_fd_sc_hd__buf_2 output509 (.A(net509),
    .X(c1_i_req_data[30]));
 sky130_fd_sc_hd__buf_2 output510 (.A(net510),
    .X(c1_i_req_data[31]));
 sky130_fd_sc_hd__buf_2 output511 (.A(net511),
    .X(c1_i_req_data[3]));
 sky130_fd_sc_hd__buf_2 output512 (.A(net512),
    .X(c1_i_req_data[4]));
 sky130_fd_sc_hd__buf_2 output513 (.A(net513),
    .X(c1_i_req_data[5]));
 sky130_fd_sc_hd__buf_2 output514 (.A(net514),
    .X(c1_i_req_data[6]));
 sky130_fd_sc_hd__buf_2 output515 (.A(net515),
    .X(c1_i_req_data[7]));
 sky130_fd_sc_hd__buf_2 output516 (.A(net516),
    .X(c1_i_req_data[8]));
 sky130_fd_sc_hd__buf_2 output517 (.A(net517),
    .X(c1_i_req_data[9]));
 sky130_fd_sc_hd__buf_2 output518 (.A(net518),
    .X(c1_i_req_data_valid));
 sky130_fd_sc_hd__buf_2 output519 (.A(net519),
    .X(c1_rst));
 sky130_fd_sc_hd__clkbuf_1 output520 (.A(net520),
    .X(dcache_clk));
 sky130_fd_sc_hd__buf_2 output521 (.A(net521),
    .X(dcache_mem_addr[0]));
 sky130_fd_sc_hd__buf_2 output522 (.A(net522),
    .X(dcache_mem_addr[10]));
 sky130_fd_sc_hd__buf_2 output523 (.A(net523),
    .X(dcache_mem_addr[11]));
 sky130_fd_sc_hd__buf_2 output524 (.A(net524),
    .X(dcache_mem_addr[12]));
 sky130_fd_sc_hd__buf_2 output525 (.A(net525),
    .X(dcache_mem_addr[13]));
 sky130_fd_sc_hd__buf_2 output526 (.A(net526),
    .X(dcache_mem_addr[14]));
 sky130_fd_sc_hd__buf_2 output527 (.A(net527),
    .X(dcache_mem_addr[15]));
 sky130_fd_sc_hd__buf_2 output528 (.A(net528),
    .X(dcache_mem_addr[16]));
 sky130_fd_sc_hd__buf_2 output529 (.A(net529),
    .X(dcache_mem_addr[17]));
 sky130_fd_sc_hd__buf_2 output530 (.A(net530),
    .X(dcache_mem_addr[18]));
 sky130_fd_sc_hd__buf_2 output531 (.A(net531),
    .X(dcache_mem_addr[19]));
 sky130_fd_sc_hd__buf_2 output532 (.A(net532),
    .X(dcache_mem_addr[1]));
 sky130_fd_sc_hd__buf_2 output533 (.A(net533),
    .X(dcache_mem_addr[20]));
 sky130_fd_sc_hd__buf_2 output534 (.A(net534),
    .X(dcache_mem_addr[21]));
 sky130_fd_sc_hd__buf_2 output535 (.A(net535),
    .X(dcache_mem_addr[22]));
 sky130_fd_sc_hd__buf_2 output536 (.A(net536),
    .X(dcache_mem_addr[23]));
 sky130_fd_sc_hd__buf_2 output537 (.A(net537),
    .X(dcache_mem_addr[2]));
 sky130_fd_sc_hd__buf_2 output538 (.A(net538),
    .X(dcache_mem_addr[3]));
 sky130_fd_sc_hd__buf_2 output539 (.A(net539),
    .X(dcache_mem_addr[4]));
 sky130_fd_sc_hd__buf_2 output540 (.A(net540),
    .X(dcache_mem_addr[5]));
 sky130_fd_sc_hd__buf_2 output541 (.A(net541),
    .X(dcache_mem_addr[6]));
 sky130_fd_sc_hd__buf_2 output542 (.A(net542),
    .X(dcache_mem_addr[7]));
 sky130_fd_sc_hd__buf_2 output543 (.A(net543),
    .X(dcache_mem_addr[8]));
 sky130_fd_sc_hd__buf_2 output544 (.A(net544),
    .X(dcache_mem_addr[9]));
 sky130_fd_sc_hd__buf_2 output545 (.A(net545),
    .X(dcache_mem_cache_enable));
 sky130_fd_sc_hd__buf_2 output546 (.A(net546),
    .X(dcache_mem_i_data[0]));
 sky130_fd_sc_hd__buf_2 output547 (.A(net547),
    .X(dcache_mem_i_data[10]));
 sky130_fd_sc_hd__buf_2 output548 (.A(net548),
    .X(dcache_mem_i_data[11]));
 sky130_fd_sc_hd__buf_2 output549 (.A(net549),
    .X(dcache_mem_i_data[12]));
 sky130_fd_sc_hd__buf_2 output550 (.A(net550),
    .X(dcache_mem_i_data[13]));
 sky130_fd_sc_hd__buf_2 output551 (.A(net551),
    .X(dcache_mem_i_data[14]));
 sky130_fd_sc_hd__buf_2 output552 (.A(net552),
    .X(dcache_mem_i_data[15]));
 sky130_fd_sc_hd__buf_2 output553 (.A(net553),
    .X(dcache_mem_i_data[1]));
 sky130_fd_sc_hd__buf_2 output554 (.A(net554),
    .X(dcache_mem_i_data[2]));
 sky130_fd_sc_hd__buf_2 output555 (.A(net555),
    .X(dcache_mem_i_data[3]));
 sky130_fd_sc_hd__buf_2 output556 (.A(net556),
    .X(dcache_mem_i_data[4]));
 sky130_fd_sc_hd__buf_2 output557 (.A(net557),
    .X(dcache_mem_i_data[5]));
 sky130_fd_sc_hd__buf_2 output558 (.A(net558),
    .X(dcache_mem_i_data[6]));
 sky130_fd_sc_hd__buf_2 output559 (.A(net559),
    .X(dcache_mem_i_data[7]));
 sky130_fd_sc_hd__buf_2 output560 (.A(net560),
    .X(dcache_mem_i_data[8]));
 sky130_fd_sc_hd__buf_2 output561 (.A(net561),
    .X(dcache_mem_i_data[9]));
 sky130_fd_sc_hd__buf_2 output562 (.A(net562),
    .X(dcache_mem_req));
 sky130_fd_sc_hd__buf_2 output563 (.A(net563),
    .X(dcache_mem_sel[0]));
 sky130_fd_sc_hd__buf_2 output564 (.A(net564),
    .X(dcache_mem_sel[1]));
 sky130_fd_sc_hd__buf_2 output565 (.A(net565),
    .X(dcache_mem_we));
 sky130_fd_sc_hd__buf_2 output566 (.A(net566),
    .X(dcache_rst));
 sky130_fd_sc_hd__buf_2 output567 (.A(net567),
    .X(dcache_wb_ack));
 sky130_fd_sc_hd__buf_2 output568 (.A(net568),
    .X(dcache_wb_err));
 sky130_fd_sc_hd__buf_2 output569 (.A(net569),
    .X(dcache_wb_i_dat[0]));
 sky130_fd_sc_hd__buf_2 output570 (.A(net570),
    .X(dcache_wb_i_dat[10]));
 sky130_fd_sc_hd__buf_2 output571 (.A(net571),
    .X(dcache_wb_i_dat[11]));
 sky130_fd_sc_hd__buf_2 output572 (.A(net572),
    .X(dcache_wb_i_dat[12]));
 sky130_fd_sc_hd__buf_2 output573 (.A(net573),
    .X(dcache_wb_i_dat[13]));
 sky130_fd_sc_hd__buf_2 output574 (.A(net574),
    .X(dcache_wb_i_dat[14]));
 sky130_fd_sc_hd__buf_2 output575 (.A(net575),
    .X(dcache_wb_i_dat[15]));
 sky130_fd_sc_hd__buf_2 output576 (.A(net576),
    .X(dcache_wb_i_dat[1]));
 sky130_fd_sc_hd__buf_2 output577 (.A(net577),
    .X(dcache_wb_i_dat[2]));
 sky130_fd_sc_hd__buf_2 output578 (.A(net578),
    .X(dcache_wb_i_dat[3]));
 sky130_fd_sc_hd__buf_2 output579 (.A(net579),
    .X(dcache_wb_i_dat[4]));
 sky130_fd_sc_hd__buf_2 output580 (.A(net580),
    .X(dcache_wb_i_dat[5]));
 sky130_fd_sc_hd__buf_2 output581 (.A(net581),
    .X(dcache_wb_i_dat[6]));
 sky130_fd_sc_hd__buf_2 output582 (.A(net582),
    .X(dcache_wb_i_dat[7]));
 sky130_fd_sc_hd__buf_2 output583 (.A(net583),
    .X(dcache_wb_i_dat[8]));
 sky130_fd_sc_hd__buf_2 output584 (.A(net584),
    .X(dcache_wb_i_dat[9]));
 sky130_fd_sc_hd__clkbuf_1 output585 (.A(net585),
    .X(ic0_clk));
 sky130_fd_sc_hd__buf_2 output586 (.A(net586),
    .X(ic0_mem_addr[0]));
 sky130_fd_sc_hd__buf_2 output587 (.A(net587),
    .X(ic0_mem_addr[10]));
 sky130_fd_sc_hd__buf_2 output588 (.A(net588),
    .X(ic0_mem_addr[11]));
 sky130_fd_sc_hd__buf_2 output589 (.A(net589),
    .X(ic0_mem_addr[12]));
 sky130_fd_sc_hd__buf_2 output590 (.A(net590),
    .X(ic0_mem_addr[13]));
 sky130_fd_sc_hd__buf_2 output591 (.A(net591),
    .X(ic0_mem_addr[14]));
 sky130_fd_sc_hd__buf_2 output592 (.A(net592),
    .X(ic0_mem_addr[15]));
 sky130_fd_sc_hd__buf_2 output593 (.A(net593),
    .X(ic0_mem_addr[1]));
 sky130_fd_sc_hd__buf_2 output594 (.A(net594),
    .X(ic0_mem_addr[2]));
 sky130_fd_sc_hd__buf_2 output595 (.A(net595),
    .X(ic0_mem_addr[3]));
 sky130_fd_sc_hd__buf_2 output596 (.A(net596),
    .X(ic0_mem_addr[4]));
 sky130_fd_sc_hd__buf_2 output597 (.A(net597),
    .X(ic0_mem_addr[5]));
 sky130_fd_sc_hd__buf_2 output598 (.A(net598),
    .X(ic0_mem_addr[6]));
 sky130_fd_sc_hd__buf_2 output599 (.A(net599),
    .X(ic0_mem_addr[7]));
 sky130_fd_sc_hd__buf_2 output600 (.A(net600),
    .X(ic0_mem_addr[8]));
 sky130_fd_sc_hd__buf_2 output601 (.A(net601),
    .X(ic0_mem_addr[9]));
 sky130_fd_sc_hd__buf_2 output602 (.A(net602),
    .X(ic0_mem_cache_flush));
 sky130_fd_sc_hd__buf_2 output603 (.A(net603),
    .X(ic0_mem_ppl_submit));
 sky130_fd_sc_hd__buf_2 output604 (.A(net604),
    .X(ic0_mem_req));
 sky130_fd_sc_hd__buf_2 output605 (.A(net605),
    .X(ic0_rst));
 sky130_fd_sc_hd__buf_2 output606 (.A(net606),
    .X(ic0_wb_ack));
 sky130_fd_sc_hd__buf_2 output607 (.A(net607),
    .X(ic0_wb_err));
 sky130_fd_sc_hd__buf_2 output608 (.A(net608),
    .X(ic0_wb_i_dat[0]));
 sky130_fd_sc_hd__buf_2 output609 (.A(net609),
    .X(ic0_wb_i_dat[10]));
 sky130_fd_sc_hd__buf_2 output610 (.A(net610),
    .X(ic0_wb_i_dat[11]));
 sky130_fd_sc_hd__buf_2 output611 (.A(net611),
    .X(ic0_wb_i_dat[12]));
 sky130_fd_sc_hd__buf_2 output612 (.A(net612),
    .X(ic0_wb_i_dat[13]));
 sky130_fd_sc_hd__buf_2 output613 (.A(net613),
    .X(ic0_wb_i_dat[14]));
 sky130_fd_sc_hd__buf_2 output614 (.A(net614),
    .X(ic0_wb_i_dat[15]));
 sky130_fd_sc_hd__buf_2 output615 (.A(net615),
    .X(ic0_wb_i_dat[1]));
 sky130_fd_sc_hd__buf_2 output616 (.A(net616),
    .X(ic0_wb_i_dat[2]));
 sky130_fd_sc_hd__buf_2 output617 (.A(net617),
    .X(ic0_wb_i_dat[3]));
 sky130_fd_sc_hd__buf_2 output618 (.A(net618),
    .X(ic0_wb_i_dat[4]));
 sky130_fd_sc_hd__buf_2 output619 (.A(net619),
    .X(ic0_wb_i_dat[5]));
 sky130_fd_sc_hd__buf_2 output620 (.A(net620),
    .X(ic0_wb_i_dat[6]));
 sky130_fd_sc_hd__buf_2 output621 (.A(net621),
    .X(ic0_wb_i_dat[7]));
 sky130_fd_sc_hd__buf_2 output622 (.A(net622),
    .X(ic0_wb_i_dat[8]));
 sky130_fd_sc_hd__buf_2 output623 (.A(net623),
    .X(ic0_wb_i_dat[9]));
 sky130_fd_sc_hd__clkbuf_1 output624 (.A(net624),
    .X(ic1_clk));
 sky130_fd_sc_hd__buf_2 output625 (.A(net625),
    .X(ic1_mem_addr[0]));
 sky130_fd_sc_hd__buf_2 output626 (.A(net626),
    .X(ic1_mem_addr[10]));
 sky130_fd_sc_hd__buf_2 output627 (.A(net627),
    .X(ic1_mem_addr[11]));
 sky130_fd_sc_hd__buf_2 output628 (.A(net628),
    .X(ic1_mem_addr[12]));
 sky130_fd_sc_hd__buf_2 output629 (.A(net629),
    .X(ic1_mem_addr[13]));
 sky130_fd_sc_hd__buf_2 output630 (.A(net630),
    .X(ic1_mem_addr[14]));
 sky130_fd_sc_hd__buf_2 output631 (.A(net631),
    .X(ic1_mem_addr[15]));
 sky130_fd_sc_hd__buf_2 output632 (.A(net632),
    .X(ic1_mem_addr[1]));
 sky130_fd_sc_hd__buf_2 output633 (.A(net633),
    .X(ic1_mem_addr[2]));
 sky130_fd_sc_hd__buf_2 output634 (.A(net634),
    .X(ic1_mem_addr[3]));
 sky130_fd_sc_hd__buf_2 output635 (.A(net635),
    .X(ic1_mem_addr[4]));
 sky130_fd_sc_hd__buf_2 output636 (.A(net636),
    .X(ic1_mem_addr[5]));
 sky130_fd_sc_hd__buf_2 output637 (.A(net637),
    .X(ic1_mem_addr[6]));
 sky130_fd_sc_hd__buf_2 output638 (.A(net638),
    .X(ic1_mem_addr[7]));
 sky130_fd_sc_hd__buf_2 output639 (.A(net639),
    .X(ic1_mem_addr[8]));
 sky130_fd_sc_hd__buf_2 output640 (.A(net640),
    .X(ic1_mem_addr[9]));
 sky130_fd_sc_hd__buf_2 output641 (.A(net641),
    .X(ic1_mem_cache_flush));
 sky130_fd_sc_hd__buf_2 output642 (.A(net642),
    .X(ic1_mem_ppl_submit));
 sky130_fd_sc_hd__buf_2 output643 (.A(net643),
    .X(ic1_mem_req));
 sky130_fd_sc_hd__buf_2 output644 (.A(net644),
    .X(ic1_rst));
 sky130_fd_sc_hd__buf_2 output645 (.A(net645),
    .X(ic1_wb_ack));
 sky130_fd_sc_hd__buf_2 output646 (.A(net646),
    .X(ic1_wb_err));
 sky130_fd_sc_hd__buf_2 output647 (.A(net647),
    .X(ic1_wb_i_dat[0]));
 sky130_fd_sc_hd__buf_2 output648 (.A(net648),
    .X(ic1_wb_i_dat[10]));
 sky130_fd_sc_hd__buf_2 output649 (.A(net649),
    .X(ic1_wb_i_dat[11]));
 sky130_fd_sc_hd__buf_2 output650 (.A(net650),
    .X(ic1_wb_i_dat[12]));
 sky130_fd_sc_hd__buf_2 output651 (.A(net651),
    .X(ic1_wb_i_dat[13]));
 sky130_fd_sc_hd__buf_2 output652 (.A(net652),
    .X(ic1_wb_i_dat[14]));
 sky130_fd_sc_hd__buf_2 output653 (.A(net653),
    .X(ic1_wb_i_dat[15]));
 sky130_fd_sc_hd__buf_2 output654 (.A(net654),
    .X(ic1_wb_i_dat[1]));
 sky130_fd_sc_hd__buf_2 output655 (.A(net655),
    .X(ic1_wb_i_dat[2]));
 sky130_fd_sc_hd__buf_2 output656 (.A(net656),
    .X(ic1_wb_i_dat[3]));
 sky130_fd_sc_hd__buf_2 output657 (.A(net657),
    .X(ic1_wb_i_dat[4]));
 sky130_fd_sc_hd__buf_2 output658 (.A(net658),
    .X(ic1_wb_i_dat[5]));
 sky130_fd_sc_hd__buf_2 output659 (.A(net659),
    .X(ic1_wb_i_dat[6]));
 sky130_fd_sc_hd__buf_2 output660 (.A(net660),
    .X(ic1_wb_i_dat[7]));
 sky130_fd_sc_hd__buf_2 output661 (.A(net661),
    .X(ic1_wb_i_dat[8]));
 sky130_fd_sc_hd__buf_2 output662 (.A(net662),
    .X(ic1_wb_i_dat[9]));
 sky130_fd_sc_hd__buf_2 output663 (.A(net663),
    .X(inner_wb_4_burst));
 sky130_fd_sc_hd__buf_2 output664 (.A(net664),
    .X(inner_wb_8_burst));
 sky130_fd_sc_hd__buf_2 output665 (.A(net665),
    .X(inner_wb_adr[0]));
 sky130_fd_sc_hd__buf_2 output666 (.A(net666),
    .X(inner_wb_adr[10]));
 sky130_fd_sc_hd__buf_2 output667 (.A(net667),
    .X(inner_wb_adr[11]));
 sky130_fd_sc_hd__buf_2 output668 (.A(net668),
    .X(inner_wb_adr[12]));
 sky130_fd_sc_hd__buf_2 output669 (.A(net669),
    .X(inner_wb_adr[13]));
 sky130_fd_sc_hd__buf_2 output670 (.A(net670),
    .X(inner_wb_adr[14]));
 sky130_fd_sc_hd__buf_2 output671 (.A(net671),
    .X(inner_wb_adr[15]));
 sky130_fd_sc_hd__buf_2 output672 (.A(net672),
    .X(inner_wb_adr[16]));
 sky130_fd_sc_hd__buf_2 output673 (.A(net673),
    .X(inner_wb_adr[17]));
 sky130_fd_sc_hd__buf_2 output674 (.A(net674),
    .X(inner_wb_adr[18]));
 sky130_fd_sc_hd__buf_2 output675 (.A(net675),
    .X(inner_wb_adr[19]));
 sky130_fd_sc_hd__buf_2 output676 (.A(net676),
    .X(inner_wb_adr[1]));
 sky130_fd_sc_hd__buf_2 output677 (.A(net677),
    .X(inner_wb_adr[20]));
 sky130_fd_sc_hd__buf_2 output678 (.A(net678),
    .X(inner_wb_adr[21]));
 sky130_fd_sc_hd__buf_2 output679 (.A(net679),
    .X(inner_wb_adr[22]));
 sky130_fd_sc_hd__buf_2 output680 (.A(net680),
    .X(inner_wb_adr[23]));
 sky130_fd_sc_hd__buf_2 output681 (.A(net681),
    .X(inner_wb_adr[2]));
 sky130_fd_sc_hd__buf_2 output682 (.A(net682),
    .X(inner_wb_adr[3]));
 sky130_fd_sc_hd__buf_2 output683 (.A(net683),
    .X(inner_wb_adr[4]));
 sky130_fd_sc_hd__buf_2 output684 (.A(net684),
    .X(inner_wb_adr[5]));
 sky130_fd_sc_hd__buf_2 output685 (.A(net685),
    .X(inner_wb_adr[6]));
 sky130_fd_sc_hd__buf_2 output686 (.A(net686),
    .X(inner_wb_adr[7]));
 sky130_fd_sc_hd__buf_2 output687 (.A(net687),
    .X(inner_wb_adr[8]));
 sky130_fd_sc_hd__buf_2 output688 (.A(net688),
    .X(inner_wb_adr[9]));
 sky130_fd_sc_hd__buf_2 output689 (.A(net689),
    .X(inner_wb_cyc));
 sky130_fd_sc_hd__buf_2 output690 (.A(net690),
    .X(inner_wb_o_dat[0]));
 sky130_fd_sc_hd__buf_2 output691 (.A(net691),
    .X(inner_wb_o_dat[10]));
 sky130_fd_sc_hd__buf_2 output692 (.A(net692),
    .X(inner_wb_o_dat[11]));
 sky130_fd_sc_hd__buf_2 output693 (.A(net693),
    .X(inner_wb_o_dat[12]));
 sky130_fd_sc_hd__buf_2 output694 (.A(net694),
    .X(inner_wb_o_dat[13]));
 sky130_fd_sc_hd__buf_2 output695 (.A(net695),
    .X(inner_wb_o_dat[14]));
 sky130_fd_sc_hd__buf_2 output696 (.A(net696),
    .X(inner_wb_o_dat[15]));
 sky130_fd_sc_hd__buf_2 output697 (.A(net697),
    .X(inner_wb_o_dat[1]));
 sky130_fd_sc_hd__buf_2 output698 (.A(net698),
    .X(inner_wb_o_dat[2]));
 sky130_fd_sc_hd__buf_2 output699 (.A(net699),
    .X(inner_wb_o_dat[3]));
 sky130_fd_sc_hd__buf_2 output700 (.A(net700),
    .X(inner_wb_o_dat[4]));
 sky130_fd_sc_hd__buf_2 output701 (.A(net701),
    .X(inner_wb_o_dat[5]));
 sky130_fd_sc_hd__buf_2 output702 (.A(net702),
    .X(inner_wb_o_dat[6]));
 sky130_fd_sc_hd__buf_2 output703 (.A(net703),
    .X(inner_wb_o_dat[7]));
 sky130_fd_sc_hd__buf_2 output704 (.A(net704),
    .X(inner_wb_o_dat[8]));
 sky130_fd_sc_hd__buf_2 output705 (.A(net705),
    .X(inner_wb_o_dat[9]));
 sky130_fd_sc_hd__buf_2 output706 (.A(net706),
    .X(inner_wb_sel[0]));
 sky130_fd_sc_hd__buf_2 output707 (.A(net707),
    .X(inner_wb_sel[1]));
 sky130_fd_sc_hd__buf_2 output708 (.A(net708),
    .X(inner_wb_stb));
 sky130_fd_sc_hd__buf_2 output709 (.A(net709),
    .X(inner_wb_we));
 sky130_fd_sc_hd__clkbuf_16 fanout710 (.A(net211),
    .X(net710));
 sky130_fd_sc_hd__conb_1 interconnect_inner_711 (.LO(net711));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_core_clock (.A(clknet_3_1_0_core_clock),
    .X(clknet_leaf_1_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_core_clock (.A(clknet_3_1_0_core_clock),
    .X(clknet_leaf_2_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_core_clock (.A(clknet_3_1_0_core_clock),
    .X(clknet_leaf_3_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_core_clock (.A(clknet_3_1_0_core_clock),
    .X(clknet_leaf_4_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_core_clock (.A(clknet_3_1_0_core_clock),
    .X(clknet_leaf_5_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_core_clock (.A(clknet_3_1_0_core_clock),
    .X(clknet_leaf_6_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_core_clock (.A(clknet_3_1_0_core_clock),
    .X(clknet_leaf_7_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_core_clock (.A(clknet_3_1_0_core_clock),
    .X(clknet_leaf_8_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_core_clock (.A(clknet_3_1_0_core_clock),
    .X(clknet_leaf_9_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_core_clock (.A(clknet_3_1_0_core_clock),
    .X(clknet_leaf_10_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_core_clock (.A(clknet_3_4_0_core_clock),
    .X(clknet_leaf_11_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_core_clock (.A(clknet_3_4_0_core_clock),
    .X(clknet_leaf_12_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_core_clock (.A(clknet_3_4_0_core_clock),
    .X(clknet_leaf_13_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_core_clock (.A(clknet_3_4_0_core_clock),
    .X(clknet_leaf_14_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_core_clock (.A(clknet_3_4_0_core_clock),
    .X(clknet_leaf_15_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_core_clock (.A(clknet_3_4_0_core_clock),
    .X(clknet_leaf_16_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_core_clock (.A(clknet_3_4_0_core_clock),
    .X(clknet_leaf_17_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_core_clock (.A(clknet_3_4_0_core_clock),
    .X(clknet_leaf_18_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_core_clock (.A(clknet_3_4_0_core_clock),
    .X(clknet_leaf_19_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_core_clock (.A(clknet_3_4_0_core_clock),
    .X(clknet_leaf_20_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_core_clock (.A(clknet_3_5_0_core_clock),
    .X(clknet_leaf_21_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_core_clock (.A(clknet_3_5_0_core_clock),
    .X(clknet_leaf_22_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_core_clock (.A(clknet_3_5_0_core_clock),
    .X(clknet_leaf_23_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_core_clock (.A(clknet_3_5_0_core_clock),
    .X(clknet_leaf_24_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_core_clock (.A(clknet_3_5_0_core_clock),
    .X(clknet_leaf_25_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_core_clock (.A(clknet_3_5_0_core_clock),
    .X(clknet_leaf_26_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_core_clock (.A(clknet_3_5_0_core_clock),
    .X(clknet_leaf_27_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_core_clock (.A(clknet_3_5_0_core_clock),
    .X(clknet_leaf_28_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_core_clock (.A(clknet_3_5_0_core_clock),
    .X(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_30_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_31_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_32_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_33_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_core_clock (.A(clknet_3_4_0_core_clock),
    .X(clknet_leaf_34_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_core_clock (.A(clknet_3_4_0_core_clock),
    .X(clknet_leaf_35_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_core_clock (.A(clknet_3_6_0_core_clock),
    .X(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_core_clock (.A(clknet_3_6_0_core_clock),
    .X(clknet_leaf_37_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_core_clock (.A(clknet_3_6_0_core_clock),
    .X(clknet_leaf_38_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_core_clock (.A(clknet_3_6_0_core_clock),
    .X(clknet_leaf_39_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_core_clock (.A(clknet_3_6_0_core_clock),
    .X(clknet_leaf_40_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_core_clock (.A(clknet_3_6_0_core_clock),
    .X(clknet_leaf_41_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_44_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_46_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_47_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_48_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_core_clock (.A(clknet_3_7_0_core_clock),
    .X(clknet_leaf_50_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_core_clock (.A(clknet_3_6_0_core_clock),
    .X(clknet_leaf_51_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_core_clock (.A(clknet_3_6_0_core_clock),
    .X(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_core_clock (.A(clknet_3_6_0_core_clock),
    .X(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_core_clock (.A(clknet_3_6_0_core_clock),
    .X(clknet_leaf_55_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_core_clock (.A(clknet_3_6_0_core_clock),
    .X(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_57_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_58_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_59_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_60_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_61_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_63_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_core_clock (.A(clknet_3_2_0_core_clock),
    .X(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_core_clock (.A(clknet_3_2_0_core_clock),
    .X(clknet_leaf_67_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_core_clock (.A(clknet_3_2_0_core_clock),
    .X(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_core_clock (.A(clknet_3_2_0_core_clock),
    .X(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_core_clock (.A(clknet_3_2_0_core_clock),
    .X(clknet_leaf_70_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_core_clock (.A(clknet_3_2_0_core_clock),
    .X(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_core_clock (.A(clknet_3_2_0_core_clock),
    .X(clknet_leaf_72_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_core_clock (.A(clknet_3_2_0_core_clock),
    .X(clknet_leaf_73_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_74_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_75_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_76_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_77_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_78_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_core_clock (.A(clknet_3_3_0_core_clock),
    .X(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_core_clock (.A(clknet_3_1_0_core_clock),
    .X(clknet_leaf_80_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_81_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_83_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_84_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_85_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_86_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_87_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_88_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_89_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_90_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_91_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_92_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_core_clock (.A(clknet_3_0_0_core_clock),
    .X(clknet_leaf_93_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_core_clock (.A(core_clock),
    .X(clknet_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_core_clock (.A(clknet_0_core_clock),
    .X(clknet_1_0_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_core_clock (.A(clknet_1_0_0_core_clock),
    .X(clknet_1_0_1_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_core_clock (.A(clknet_0_core_clock),
    .X(clknet_1_1_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_core_clock (.A(clknet_1_1_0_core_clock),
    .X(clknet_1_1_1_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_core_clock (.A(clknet_1_0_1_core_clock),
    .X(clknet_2_0_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_core_clock (.A(clknet_1_0_1_core_clock),
    .X(clknet_2_1_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_core_clock (.A(clknet_1_1_1_core_clock),
    .X(clknet_2_2_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_core_clock (.A(clknet_1_1_1_core_clock),
    .X(clknet_2_3_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_core_clock (.A(clknet_2_0_0_core_clock),
    .X(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_core_clock (.A(clknet_2_0_0_core_clock),
    .X(clknet_3_1_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_core_clock (.A(clknet_2_1_0_core_clock),
    .X(clknet_3_2_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_core_clock (.A(clknet_2_1_0_core_clock),
    .X(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_core_clock (.A(clknet_2_2_0_core_clock),
    .X(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_core_clock (.A(clknet_2_2_0_core_clock),
    .X(clknet_3_5_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_core_clock (.A(clknet_2_3_0_core_clock),
    .X(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_core_clock (.A(clknet_2_3_0_core_clock),
    .X(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_core_clock (.A(clknet_3_2_0_core_clock),
    .X(clknet_opt_1_0_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_core_clock (.A(clknet_3_6_0_core_clock),
    .X(clknet_opt_2_0_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_1_core_clock (.A(clknet_opt_2_0_core_clock),
    .X(clknet_opt_2_1_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__A3 (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__B (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__B (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A2 (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__C1 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__C1 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__C1 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__C1 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__A (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__A (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__A (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__C1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__C1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__B (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__B (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__S (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3228__A (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__A (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__A (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__C (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__B2 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__B1 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__A1 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__B1 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__B2 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__B (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__B (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__B (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__B (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__A (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__B (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__B (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__B (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__B (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__B (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__B (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__B (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__B (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__B (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__B (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__A (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3223__A (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__A (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__B (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__B (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__S (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__B1 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__B1 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__C1 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__B1 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__B1 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__B (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__B (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__A (.DIODE(_0836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__A (.DIODE(_0837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A (.DIODE(_0838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A (.DIODE(_0838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A (.DIODE(_0838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__A (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__S (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__S (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__S (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__S (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__S (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__A (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__B (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__B1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3376__B1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__B1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__S (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__S (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__S (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__S (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__S (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__S (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__A (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__A (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__A (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__A (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__S (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__S (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__S (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__S (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__S (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__S (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__S (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__S (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__S (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__S (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__A (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__A (.DIODE(_0849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__A (.DIODE(_0851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__A (.DIODE(_0852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__A (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__C1 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A1 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__C1 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__B1 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__B1 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__B1 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__B1 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__S (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__C1 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3262__A (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__C1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__C1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__A (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3411__A (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__S (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__S (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__B1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__C1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__A1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__A1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__S (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__S (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__S (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__S (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__S (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__S (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__S (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__A (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__S (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__A (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__S (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__S (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__S (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__S (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__S (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__S (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__S (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__A (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__A (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__A (.DIODE(_0857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__S (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__S (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__S0 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__S1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__A (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__A1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__A (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__S1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__A (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__A (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__S1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__S1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__S1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__S1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__S1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__S1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__S1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__S1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__S1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__S1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__S1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__S1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__S1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__S1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__S1 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__S1 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__S1 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__S1 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__S1 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__S1 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__S1 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__A0 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__A (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__A (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__S0 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__S (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__S (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__S0 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__S0 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__S (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__S0 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__S (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3289__S (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__S (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A1 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A1 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__A1 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A1 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A1 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__A (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__A1 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3276__A (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A1 (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__A (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A1 (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A1 (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__A1 (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__A1 (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__A1 (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__A (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__A1 (.DIODE(_0869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__A1 (.DIODE(_0872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A1 (.DIODE(_0872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__B1 (.DIODE(_0872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__B1 (.DIODE(_0872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__B1 (.DIODE(_0872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__S (.DIODE(_0872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__A (.DIODE(_0872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__A1 (.DIODE(_0872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__A (.DIODE(_0872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__B1 (.DIODE(_0872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__C1 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__C1 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__B1 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__C1 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A1 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__C1 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__B1 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__A1 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__B1 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__C1 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__B2 (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__S (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__S (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__S (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A1 (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__A1 (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__A1 (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3376__A1 (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__A1 (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A1 (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__S (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__C1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__A1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__S (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__S (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__A1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__S (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__S0 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__S0 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__S0 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__S0 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__S0 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__S0 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__S0 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__S0 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__A (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__S0 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__S0 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__S0 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__S0 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__S0 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__S0 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__S0 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__S0 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__S0 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__A1 (.DIODE(_0892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__A2 (.DIODE(_0894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__S0 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__S (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__S (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__S (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__S (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__S0 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__S0 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__S (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__S (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__A (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__S (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__S (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__S (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__S0 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__S0 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__S0 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__S0 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__S (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__A (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__A (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__S0 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__S0 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__S0 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__S0 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__S0 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__S0 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__S0 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__S0 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__S0 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__S (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__S0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__S0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__S0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__S0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__S0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__S0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__S0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__S0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__A0 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__S0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__S0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__S0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__S0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__S (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__S (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__S (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__A (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__S0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__S0 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__A1 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__A1 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__S1 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__A (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__A (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__S1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__S1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__S1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__S1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__S1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__S1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__S1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__S1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__S1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__S1 (.DIODE(_0902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A1 (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A1 (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__B1 (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__C1 (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__C1 (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__C1 (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__A1 (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__B1 (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__B1 (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__A (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__C1 (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__C1 (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__S (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__A (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__S (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__S (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__B1 (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__A1 (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__C1 (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__S (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A1 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A1 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__A1 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A1 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__A1 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__A (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A1 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3316__A (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A1 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__A1 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A1 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A1 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A1 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__A1 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3360__A (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__A1 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__S0 (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__S0 (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__S0 (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__S (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__A (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__S1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__S1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__S1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__S1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__S1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__S1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__A (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__S1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__S1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__S1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__S1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__S1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__S1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__C1 (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__C1 (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__C1 (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__A1 (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__B1 (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__S (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__S (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__S (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__A (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__S (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__S (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__S (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__C1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__A1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__A1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__C1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__S (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__A1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__C1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__B2 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__A1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__A1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__C (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__B1 (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__A1 (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__A1 (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__B1 (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__A2 (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A2 (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__S (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__A1 (.DIODE(_0943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__A2 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__A2 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__A (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__A (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__S1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__S1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__S1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__S1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__S1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__S1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__A1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__S1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A1 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__B2 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__B2 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__C1 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__B1 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__B1 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__C1 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__B2 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__A1 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__A (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A1 (.DIODE(_0963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A2 (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__A1 (.DIODE(_0980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__A2 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A2 (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__B (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__B (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__B (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__B (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__B (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__B (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__B (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A1 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A1 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A1 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__B1 (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A2 (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A3 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__B1 (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__B1 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__C1 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__B2 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A2 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__C1 (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__B (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__A1_N (.DIODE(_1065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__A2_N (.DIODE(_1069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__A0 (.DIODE(_1072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__B1 (.DIODE(_1078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__B (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A1 (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A1 (.DIODE(_1088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A2 (.DIODE(_1088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A3 (.DIODE(_1095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A2 (.DIODE(_1098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__B (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A2 (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A2 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A2 (.DIODE(_1137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__B (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__S0 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__S0 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A2 (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A3 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__B (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A2 (.DIODE(_1168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__S (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__S (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__S (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__S (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__S (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__S (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__S (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__S (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__S (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__S (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__A2 (.DIODE(_1178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__B (.DIODE(_1179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__A3 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A2 (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__A0 (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__C (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A0 (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__B1 (.DIODE(_1220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__B (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__B (.DIODE(_1268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__C_N (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__D (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__A1 (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__B1 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__A1 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__S (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__S (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__S (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__S (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__S (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__S (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__S (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__S (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__S (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__S (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A (.DIODE(_1325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A (.DIODE(_1336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__B (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__B (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__B (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__B (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__B (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__B (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__B (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__B1 (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__C1 (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__B1 (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__C1 (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__B1 (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__S (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__S (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__S (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__S (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__S (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A1 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__A (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__A (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A1 (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__A (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A1 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A1 (.DIODE(_1385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A (.DIODE(_1387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A1 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__S (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__S (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__S (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__S (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__S (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__S (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__S (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__S (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__S (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__S (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A1 (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A (.DIODE(_1392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A1 (.DIODE(_1395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__A1 (.DIODE(_1397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A1 (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A1 (.DIODE(_1405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__S0 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__S0 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__S (.DIODE(_1408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__S (.DIODE(_1408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__S (.DIODE(_1408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__S (.DIODE(_1408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__A (.DIODE(_1408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__S (.DIODE(_1408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__S (.DIODE(_1408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__S (.DIODE(_1408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__S (.DIODE(_1408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A (.DIODE(_1408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__S (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__S (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__S0 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__S0 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__S0 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__S0 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__S0 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__S0 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__S0 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__A (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__B1 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__A1 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__B (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__B (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__C_N (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__A (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__C (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__B2 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__B2 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__A1 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A1 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A1 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__A1 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__B1 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__C1 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__B (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A0 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__C1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__C1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__C1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__B1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__B (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__B1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__S (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__A (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__A1 (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__A1 (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__S1 (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A1 (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__S1 (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__A1 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__A (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__A (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__S1 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__S1 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__S1 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__S1 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__S1 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A1 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__A (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__A1 (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__A1 (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__A (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__A (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__A1 (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A1 (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__A (.DIODE(_1423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A1 (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__A (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__A (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__A (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__A1 (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A1 (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A1 (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__A1 (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__A2 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__A (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__A (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__A1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__A1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__S1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__S1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A1 (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__A1 (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__B1 (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__C1 (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__C1 (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__C1 (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__B1 (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__C1 (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__B1 (.DIODE(_1432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A3 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__S (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__S (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__S (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__S (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__S0 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__S0 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__S0 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__S0 (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A (.DIODE(_1437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__S (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__S (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__S (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__S (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__S (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__S (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__S (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__S0 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__S0 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__S0 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__S (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__S0 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A1 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A1 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__B2 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__C1 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__C1 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__B1 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A2 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A1 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__S1 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__S1 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__S (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__S (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__S (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__S (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__S (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__S (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__S (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__S (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__S (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__A (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__A (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4149__A (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__B2 (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__B2 (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__A1 (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__S (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__S (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__S (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A1 (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__B_N (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__S (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__A (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__A1 (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__B_N (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__S (.DIODE(_1448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__C1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__C1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__C1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__C1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__B1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__C1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__B1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__S (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__S (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__S (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__S (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__S (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__S (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__S0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__S0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__S0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__S0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A1 (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__A1 (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__A (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__S1 (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__S1 (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__B1 (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__S1 (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__S1 (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__S1 (.DIODE(_1454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__C1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__C1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__B2 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__B1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__C1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__B2 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__C1 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A1 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__A (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__C1 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__C1 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__A1 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__C1 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A1 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__C1 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A1 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A2 (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__A (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__B2 (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A1 (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__B1 (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__B1 (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__B1 (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__B1 (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__B1 (.DIODE(_1464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A2 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__S (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__S (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__S (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__S (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__S0 (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__S (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__S (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__S (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__S0 (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A2 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A2 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A1 (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__A (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__A1 (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__A1 (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__A (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__A (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A1 (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__C1 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__A1 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__C1 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A1 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__A1 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A1 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A1 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__S0 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__B1 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A1 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__S0 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__S0 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A3 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__C (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__S0 (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__S0 (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A2 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__A (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__A (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__S1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__A1 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__B2 (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__B1 (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A2 (.DIODE(_1505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A2 (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A2 (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A2 (.DIODE(_1510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__B1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A3 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__B1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__C1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__C1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__A1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__B1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__B1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__C1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__A1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__B1 (.DIODE(_1521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__A1 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A1 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__A (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A1 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__A1 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A1 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__A1 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A1 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__S (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__S (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__S (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4310__S (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__S (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__S (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__S (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__S (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__S (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__S (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__B1 (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__C1 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__B1 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__A1 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__C1 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__B1 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__C1 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__B2 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A1 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A1 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__C1 (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__B1 (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A (.DIODE(_1534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__B1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__C1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__C1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__C1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__B1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__A1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__B1 (.DIODE(_1540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__A2 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__A0 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__B1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__B1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__C1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__C1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__A1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__C1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__C1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__C1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__C1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__B1 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A2 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__A1 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__A1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__A1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__A1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__S1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__S1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__S1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__S1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__A1 (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A2 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__B (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__B (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__C1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__C1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__A1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__C1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__C1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__C1 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__A (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__A (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__A1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__A1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__A1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__A (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__S1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A2 (.DIODE(_1582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__A (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__A (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A1 (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A1 (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__A1 (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__A (.DIODE(_1584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A2 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__B (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A2 (.DIODE(_1600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__S0 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__S0 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__S0 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__B1 (.DIODE(_1613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__B1 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A (.DIODE(_1619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__A2 (.DIODE(_1623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__B (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__B (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__A2 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A2 (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A2 (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__B1 (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__B1 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A2 (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__B (.DIODE(_1663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__B2 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__B1 (.DIODE(_1704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__B (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__A2 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__A2 (.DIODE(_1716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__B1 (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__B1_N (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__A2 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__B1 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__B (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__A2_N (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__A2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__A2 (.DIODE(_1791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A2 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__B (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A2 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__B1 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__B1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__B (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A3 (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__B1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__B2 (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__B1 (.DIODE(_1841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A2 (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__B1 (.DIODE(_1854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A2 (.DIODE(_1864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__A3 (.DIODE(_1880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__A1_N (.DIODE(_1885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__A2_N (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A1 (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A1 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__A (.DIODE(_1893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A1 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__A (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A (.DIODE(_1896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A (.DIODE(_1896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__A (.DIODE(_1896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__A (.DIODE(_1896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A (.DIODE(_1896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__A (.DIODE(_1897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A (.DIODE(_1897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A (.DIODE(_1897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__A (.DIODE(_1897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__A (.DIODE(_1897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A (.DIODE(_1897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A (.DIODE(_1897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A (.DIODE(_1897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__A (.DIODE(_1897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A (.DIODE(_1897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A1 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A1 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__A1 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__A1 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__A1 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A1 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A1 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__A (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__B1_N (.DIODE(_1899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__A1 (.DIODE(_1899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__B (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__A (.DIODE(_1901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__A (.DIODE(_1909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__C1 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__C1 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__C1 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__B1 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__B1 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A1 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A1 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A1 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A1 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A1 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__A (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A (.DIODE(_1921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A (.DIODE(_1921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A (.DIODE(_1921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__A (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__B (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__A3 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A3 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A3 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__A3 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A3 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A3 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A3 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A3 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A3 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A3 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__A1_N (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A1 (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__A0 (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__A (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__A (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__B (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__B (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__B (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__B (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__B (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__B (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__B (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__B (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__B (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__B (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__B (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A1 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__A (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A1 (.DIODE(_1935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A (.DIODE(_1935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A (.DIODE(_1935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A (.DIODE(_1935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A (.DIODE(_1935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A (.DIODE(_1935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A (.DIODE(_1935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__A (.DIODE(_1935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A (.DIODE(_1935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A (.DIODE(_1935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A1 (.DIODE(_1937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A (.DIODE(_1937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A (.DIODE(_1937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A (.DIODE(_1937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A (.DIODE(_1937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A (.DIODE(_1937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A (.DIODE(_1937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__A (.DIODE(_1937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A (.DIODE(_1937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__A (.DIODE(_1937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__A1 (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A1 (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A1 (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__A1 (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A1 (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__A1 (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A1 (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A1 (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__A1 (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A1 (.DIODE(_1939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A1 (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A (.DIODE(_1940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A1 (.DIODE(_1942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A (.DIODE(_1942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A (.DIODE(_1942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A (.DIODE(_1942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A (.DIODE(_1942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A (.DIODE(_1942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A (.DIODE(_1942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A (.DIODE(_1942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A (.DIODE(_1942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A (.DIODE(_1942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A1 (.DIODE(_1944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A (.DIODE(_1944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A (.DIODE(_1944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A (.DIODE(_1944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A (.DIODE(_1944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A (.DIODE(_1944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A (.DIODE(_1944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__A (.DIODE(_1944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A (.DIODE(_1944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A (.DIODE(_1944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A1 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A1 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A1 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A1 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A1 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A1 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A1 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A1 (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__A (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__A (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A1 (.DIODE(_1948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A1 (.DIODE(_1948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__A1 (.DIODE(_1948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A1 (.DIODE(_1948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A1 (.DIODE(_1948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__A1 (.DIODE(_1948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A1 (.DIODE(_1948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A1 (.DIODE(_1948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__A (.DIODE(_1948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A (.DIODE(_1948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__A1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__A1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__A (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__A (.DIODE(_1958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A (.DIODE(_1958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A (.DIODE(_1958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A (.DIODE(_1958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__A (.DIODE(_1958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__A (.DIODE(_1961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A (.DIODE(_1961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__B (.DIODE(_1961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__B (.DIODE(_1961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A3 (.DIODE(_1963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A3 (.DIODE(_1963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A3 (.DIODE(_1963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__B (.DIODE(_1963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__A (.DIODE(_1963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A3 (.DIODE(_1964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__A3 (.DIODE(_1964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__A3 (.DIODE(_1964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A3 (.DIODE(_1964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__A3 (.DIODE(_1964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A3 (.DIODE(_1964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__A3 (.DIODE(_1964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A3 (.DIODE(_1964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A3 (.DIODE(_1964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__A3 (.DIODE(_1964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__A1 (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__A1 (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A1 (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__A1 (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A1 (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A1 (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A1 (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__A1 (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__A (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A (.DIODE(_1967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__B (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__B (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__B (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__B (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__B (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__B (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__B (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__B (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__B (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__B (.DIODE(_1970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A1 (.DIODE(_1972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A1 (.DIODE(_1972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A1 (.DIODE(_1972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A1 (.DIODE(_1972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A1 (.DIODE(_1972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__A1 (.DIODE(_1972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A1 (.DIODE(_1972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A1 (.DIODE(_1972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__A (.DIODE(_1972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__A (.DIODE(_1972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__A1 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A1 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A1 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A1 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A1 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A1 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A1 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__A1 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__A (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A1 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A1 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A1 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A1 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A1 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__A1 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__A1 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A1 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__A1 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A1 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__A1 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__A1 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A1 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__A1 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__A1 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__A1 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A1 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__A1 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__A (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A1 (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__A1 (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A1 (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A1 (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A1 (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A1 (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A1 (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A1 (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__A (.DIODE(_1979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__A1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__A1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__A1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__A (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__A (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__A (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A1 (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__A (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A1 (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A1 (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__A1 (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A1 (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A1 (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__A (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__A (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__A1 (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__A (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A1 (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A1 (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A1 (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A1 (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A1 (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__A (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__A (.DIODE(_1987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__A (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__A1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__A (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A (.DIODE(_1991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__A (.DIODE(_1991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A (.DIODE(_1991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A (.DIODE(_1991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A (.DIODE(_1991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A (.DIODE(_1991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__A (.DIODE(_1991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__A (.DIODE(_1991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A (.DIODE(_1991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__A (.DIODE(_1991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A1 (.DIODE(_1995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__A1 (.DIODE(_1995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A (.DIODE(_1995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A (.DIODE(_1995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A1 (.DIODE(_1995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A1 (.DIODE(_1995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A1 (.DIODE(_1995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A1 (.DIODE(_1995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__A1 (.DIODE(_1995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__A (.DIODE(_1995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__A1 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__A1 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A1 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__A1 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__A1 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__A1 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A1 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__A1 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A1 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A1 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__B (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__A (.DIODE(_1998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__A (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__A (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__A (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__A (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__A (.DIODE(_2000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A (.DIODE(_2000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__A (.DIODE(_2000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A (.DIODE(_2000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A (.DIODE(_2000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A (.DIODE(_2000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__A (.DIODE(_2000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__A (.DIODE(_2000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A (.DIODE(_2000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__B (.DIODE(_2000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__A2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__A2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__A2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__A2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A2 (.DIODE(_2002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__C (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__C (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__C (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__C (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__C (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__C (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__C (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__C (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__C (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__C (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A1 (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__A1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__A1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__A1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__A1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__A1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__A1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__A1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__A1 (.DIODE(_2008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A1 (.DIODE(_2010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__A1 (.DIODE(_2010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__A1 (.DIODE(_2010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__A1 (.DIODE(_2010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__A1 (.DIODE(_2010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__A1 (.DIODE(_2010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A1 (.DIODE(_2010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A1 (.DIODE(_2010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__A1 (.DIODE(_2010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A1 (.DIODE(_2010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A1 (.DIODE(_2012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A1 (.DIODE(_2012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A1 (.DIODE(_2012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A1 (.DIODE(_2012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A1 (.DIODE(_2012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__A1 (.DIODE(_2012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__A1 (.DIODE(_2012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__A1 (.DIODE(_2012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A1 (.DIODE(_2012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__A1 (.DIODE(_2012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A1 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A1 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__A1 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__A1 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__A1 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A1 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A1 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A1 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A1 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__A1 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A1 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A1 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A1 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A1 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A1 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A1 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A1 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__A1 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__A1 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A1 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A (.DIODE(_2017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__A (.DIODE(_2017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A (.DIODE(_2017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A (.DIODE(_2017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A (.DIODE(_2017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A (.DIODE(_2017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__A (.DIODE(_2017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A (.DIODE(_2017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A (.DIODE(_2017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A (.DIODE(_2017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__A1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__A1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__A1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A1 (.DIODE(_2019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__A1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__A1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__A1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__A1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__A1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A1 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A1 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__A1 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A1 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__A1 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A1 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__A1 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A1 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A1 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__A1 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A1 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__A1 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A1 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A1 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__A1 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A1 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A1 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A1 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A1 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A1 (.DIODE(_2025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__B (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__B (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__B (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__B (.DIODE(_2028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A2 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__A2 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__A2 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__A2 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A2 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A2 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__A2 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A2 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A2 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A2 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__C (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__C (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__C (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__C (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__C (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__C (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__C (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__C (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__C (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__C (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__A (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__A (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__A (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__A (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__A (.DIODE(_2038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__B (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__B (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__B (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__B (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A2 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__A2 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__A2 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__A2 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A2 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__A2 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A2 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__A2 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__A2 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__A2 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__C (.DIODE(_2049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__C (.DIODE(_2049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__C (.DIODE(_2049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__C (.DIODE(_2049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__C (.DIODE(_2049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__C (.DIODE(_2049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__C (.DIODE(_2049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__C (.DIODE(_2049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__C (.DIODE(_2049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__C (.DIODE(_2049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__A (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__A (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__A (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__A (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__A (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__A (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__A (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__B (.DIODE(_2064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__B (.DIODE(_2064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__B (.DIODE(_2064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__B (.DIODE(_2064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__C (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__C (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__C (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__C (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__C (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__C (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__C (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__C (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__C (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__C (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__A (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__A (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__A (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__A (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__A (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__B (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__B (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__B (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__B (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A2 (.DIODE(_2083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A2 (.DIODE(_2083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A2 (.DIODE(_2083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A2 (.DIODE(_2083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A2 (.DIODE(_2083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__A2 (.DIODE(_2083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__A2 (.DIODE(_2083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__A2 (.DIODE(_2083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__A2 (.DIODE(_2083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__A2 (.DIODE(_2083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__A (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__A (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__A (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__A (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__A (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__C (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__C (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__C (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__C (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__C (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__C (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__C (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__C (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__C (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__C (.DIODE(_2086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__A (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__A (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__A (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__A (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__A (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__A (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__A (.DIODE(_2089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__B (.DIODE(_2099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__B (.DIODE(_2099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A (.DIODE(_2099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__B (.DIODE(_2099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__B (.DIODE(_2099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__A2 (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__A2 (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__A2 (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A2 (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__A2 (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A2 (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__A2 (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__A2 (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__A2 (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__A2 (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__C (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__C (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__C (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__C (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__C (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__C (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__C (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__C (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__C (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__C (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__A (.DIODE(_2105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__A (.DIODE(_2105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A (.DIODE(_2105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A (.DIODE(_2105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__A (.DIODE(_2105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__A (.DIODE(_2105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A (.DIODE(_2105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__A (.DIODE(_2105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__A (.DIODE(_2105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__A (.DIODE(_2105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__A (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__A (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__A (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__A (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__A (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__A (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__B (.DIODE(_2118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__B (.DIODE(_2118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__B (.DIODE(_2118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__B (.DIODE(_2118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A2 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A2 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A2 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A2 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__A2 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A2 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__A2 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__A2 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__A2 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__A2 (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__A (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__A (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__A (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__A (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__C (.DIODE(_2123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__C (.DIODE(_2123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__C (.DIODE(_2123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__C (.DIODE(_2123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__C (.DIODE(_2123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__C (.DIODE(_2123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__C (.DIODE(_2123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__C (.DIODE(_2123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__C (.DIODE(_2123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__C (.DIODE(_2123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__A (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__A (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__A (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__A (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__A (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A (.DIODE(_2134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__B (.DIODE(_2136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__B (.DIODE(_2136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__B (.DIODE(_2136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__B (.DIODE(_2136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__A2 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__A2 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A2 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A2 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__A2 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A2 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__A2 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__A2 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__A2 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A2 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__C (.DIODE(_2140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__C (.DIODE(_2140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__C (.DIODE(_2140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__C (.DIODE(_2140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__C (.DIODE(_2140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__C (.DIODE(_2140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__C (.DIODE(_2140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__C (.DIODE(_2140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__C (.DIODE(_2140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__C (.DIODE(_2140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__A (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__A (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__A (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__A (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__A (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__A (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A (.DIODE(_2150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__B (.DIODE(_2153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__B (.DIODE(_2153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__B (.DIODE(_2153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__B (.DIODE(_2153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A2 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A2 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A2 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A2 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A2 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A2 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__A2 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__A2 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A2 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__A2 (.DIODE(_2155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__C (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__C (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__C (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__C (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__C (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__C (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__C (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__C (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__C (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__C (.DIODE(_2157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__A (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__A (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__A (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__A (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__B (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__B (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__B (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__B (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A2 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A2 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A2 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A2 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A2 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A2 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A2 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A2 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__A2 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__A2 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__C (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__C (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__C (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__C (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__C (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__C (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__C (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__C (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__C (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__C (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__A (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__A (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__A (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__A (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__A (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__A (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__A (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__B (.DIODE(_2187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__B (.DIODE(_2187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__B (.DIODE(_2187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A2 (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A2 (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A2 (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A2 (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A2 (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__A2 (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__A2 (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A2 (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__A2 (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__A2 (.DIODE(_2189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__A (.DIODE(_2190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A (.DIODE(_2190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__A (.DIODE(_2190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__A (.DIODE(_2190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__A (.DIODE(_2190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__A (.DIODE(_2190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A (.DIODE(_2190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A (.DIODE(_2190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A (.DIODE(_2190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A (.DIODE(_2190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__B1 (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__B1 (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__B1 (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__B1 (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__B1 (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__B1 (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__B1 (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__B1 (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__B1 (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__B1 (.DIODE(_2192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__B (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__B (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__B (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__B (.DIODE(_2193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A2 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A2 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__A2 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__A2 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A2 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A2 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A2 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A2 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A2 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A2 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__C (.DIODE(_2197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__C (.DIODE(_2197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__C (.DIODE(_2197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__C (.DIODE(_2197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__C (.DIODE(_2197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__C (.DIODE(_2197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__C (.DIODE(_2197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__C (.DIODE(_2197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__C (.DIODE(_2197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__C (.DIODE(_2197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__A (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__A (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A (.DIODE(_2204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A1 (.DIODE(_2210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A1 (.DIODE(_2210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__A1 (.DIODE(_2210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A1 (.DIODE(_2210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A1 (.DIODE(_2210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A1 (.DIODE(_2210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__A0 (.DIODE(_2210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A1 (.DIODE(_2210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A1 (.DIODE(_2210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__A (.DIODE(_2210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A1 (.DIODE(_2211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A1 (.DIODE(_2211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A1 (.DIODE(_2211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A1 (.DIODE(_2211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(_2211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A1 (.DIODE(_2211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A1 (.DIODE(_2211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A1 (.DIODE(_2211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A1 (.DIODE(_2211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A1 (.DIODE(_2211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__D (.DIODE(_2212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__B (.DIODE(_2212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A (.DIODE(_2212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A (.DIODE(_2212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__A (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__B (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__B (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A (.DIODE(_2215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__A (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__B (.DIODE(_2217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__A2 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A2 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__A2 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A2 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A2 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__A2 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A2 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A2 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A2 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A2 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__C (.DIODE(_2221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__C (.DIODE(_2221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__C (.DIODE(_2221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__C (.DIODE(_2221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__C (.DIODE(_2221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__C (.DIODE(_2221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__C (.DIODE(_2221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__C (.DIODE(_2221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__C (.DIODE(_2221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__C (.DIODE(_2221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A1 (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A1 (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__A1 (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A1 (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A1 (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A1 (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A1 (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A1 (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A1 (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A (.DIODE(_2223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A1 (.DIODE(_2224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A1 (.DIODE(_2224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A1 (.DIODE(_2224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A1 (.DIODE(_2224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A1 (.DIODE(_2224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A1 (.DIODE(_2224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A1 (.DIODE(_2224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A1 (.DIODE(_2224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A1 (.DIODE(_2224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A1 (.DIODE(_2224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__A1 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A1 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A1 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__A1 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A1 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A1 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A0 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A1 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A1 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__A1 (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A1 (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A1 (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A1 (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A1 (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A1 (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A0 (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A1 (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A1 (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__A (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A1 (.DIODE(_2230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A1 (.DIODE(_2230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A1 (.DIODE(_2230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A1 (.DIODE(_2230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A1 (.DIODE(_2230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A1 (.DIODE(_2230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A1 (.DIODE(_2230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A1 (.DIODE(_2230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A1 (.DIODE(_2230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A1 (.DIODE(_2230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A1 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A1 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A1 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A1 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A1 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A1 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A0 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__A1 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A1 (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A (.DIODE(_2232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__A1 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A1 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A1 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A1 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A1 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A1 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A1 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A1 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A1 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__A1 (.DIODE(_2233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A1 (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A1 (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A1 (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A1 (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A1 (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A1 (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A0 (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A1 (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A1 (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A (.DIODE(_2235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A1 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A1 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A1 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A1 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A1 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A1 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A1 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A1 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A1 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A1 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__A (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__A (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__A (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__A (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__A (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__A (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__A (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A (.DIODE(_2237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A1 (.DIODE(_2239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__A1 (.DIODE(_2239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A1 (.DIODE(_2239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__A1 (.DIODE(_2239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A1 (.DIODE(_2239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A1 (.DIODE(_2239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A0 (.DIODE(_2239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A1 (.DIODE(_2239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A1 (.DIODE(_2239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A (.DIODE(_2239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__A1 (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A1 (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A1 (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A1 (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A1 (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A1 (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A0 (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A1 (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A1 (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__A (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__A1 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A1 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A1 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A1 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A1 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A1 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A1 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A1 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A1 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__A1 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A1 (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A1 (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A1 (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A1 (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A1 (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A1 (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A1 (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__A1 (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A1 (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A1 (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__A1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A1 (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A1 (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A1 (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A1 (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A1 (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A1 (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A1 (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A1 (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A1 (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__A1 (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A1 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A1 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A1 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A1 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A1 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A1 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A1 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A1 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A1 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__A1 (.DIODE(_2251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A1 (.DIODE(_2253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A1 (.DIODE(_2253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A1 (.DIODE(_2253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A1 (.DIODE(_2253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A1 (.DIODE(_2253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A1 (.DIODE(_2253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A1 (.DIODE(_2253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A1 (.DIODE(_2253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A1 (.DIODE(_2253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__A1 (.DIODE(_2253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__B (.DIODE(_2255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__B (.DIODE(_2255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__B (.DIODE(_2255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__B (.DIODE(_2255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__C (.DIODE(_2259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__C (.DIODE(_2259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__C (.DIODE(_2259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__C (.DIODE(_2259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__C (.DIODE(_2259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__C (.DIODE(_2259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__C (.DIODE(_2259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__C (.DIODE(_2259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__C (.DIODE(_2259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__C (.DIODE(_2259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__A (.DIODE(_2262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A (.DIODE(_2262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__A (.DIODE(_2262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A (.DIODE(_2262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A (.DIODE(_2262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A (.DIODE(_2262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__A (.DIODE(_2262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A (.DIODE(_2262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A (.DIODE(_2262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__A (.DIODE(_2262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__B (.DIODE(_2272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__B (.DIODE(_2272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__D (.DIODE(_2272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__B (.DIODE(_2272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A2 (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A2 (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__A2 (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__A2 (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A2 (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__A2 (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A2 (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A2 (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A2 (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__A2_N (.DIODE(_2274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__B1 (.DIODE(_2277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__B1 (.DIODE(_2277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__B1 (.DIODE(_2277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__B1 (.DIODE(_2277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__B1 (.DIODE(_2277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__B1 (.DIODE(_2277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__B1 (.DIODE(_2277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__B1 (.DIODE(_2277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__B1 (.DIODE(_2277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__B1 (.DIODE(_2277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__B (.DIODE(_2278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__B (.DIODE(_2278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__B (.DIODE(_2278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__B (.DIODE(_2278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A2 (.DIODE(_2280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A2 (.DIODE(_2280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A2 (.DIODE(_2280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A2 (.DIODE(_2280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A2 (.DIODE(_2280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__A2 (.DIODE(_2280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A2 (.DIODE(_2280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A2 (.DIODE(_2280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__A2 (.DIODE(_2280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A2 (.DIODE(_2280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__C (.DIODE(_2282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__C (.DIODE(_2282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__C (.DIODE(_2282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__C (.DIODE(_2282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__C (.DIODE(_2282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__C (.DIODE(_2282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__C (.DIODE(_2282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__C (.DIODE(_2282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__C (.DIODE(_2282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__C (.DIODE(_2282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__A (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__A (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__A (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__A (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__B (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__B (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__B (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__B (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A3 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A3 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A3 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A3 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A3 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A3 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A3 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A3 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A3 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A3 (.DIODE(_2298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__A (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A1 (.DIODE(_2301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A1 (.DIODE(_2301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A1 (.DIODE(_2301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A1 (.DIODE(_2301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A1 (.DIODE(_2301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A1 (.DIODE(_2301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A1 (.DIODE(_2301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A1 (.DIODE(_2301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A1 (.DIODE(_2301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A1 (.DIODE(_2301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__B (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__B (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__B (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__B (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__B (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__B (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__B (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__B (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__B (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__A (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__A (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A (.DIODE(_2310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A (.DIODE(_2314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A (.DIODE(_2314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A (.DIODE(_2314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A (.DIODE(_2314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A (.DIODE(_2314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A (.DIODE(_2314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A (.DIODE(_2314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A (.DIODE(_2314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A (.DIODE(_2314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A (.DIODE(_2314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A1 (.DIODE(_2316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A1 (.DIODE(_2316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A1 (.DIODE(_2316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A1 (.DIODE(_2316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A1 (.DIODE(_2316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A1 (.DIODE(_2316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A1 (.DIODE(_2316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A1 (.DIODE(_2316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A1 (.DIODE(_2316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A1 (.DIODE(_2316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__B (.DIODE(_2318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__B (.DIODE(_2318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__B (.DIODE(_2318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__B (.DIODE(_2318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A3 (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A3 (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A3 (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A3 (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A3 (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A3 (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A3 (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A3 (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A3 (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A3 (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__B (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__B (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__B (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__B (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__B (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__B (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__B (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__B (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__B (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__B (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__B (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__B (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__B (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__B (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A3 (.DIODE(_2336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A3 (.DIODE(_2336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A3 (.DIODE(_2336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A3 (.DIODE(_2336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A3 (.DIODE(_2336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A3 (.DIODE(_2336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A3 (.DIODE(_2336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A3 (.DIODE(_2336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A3 (.DIODE(_2336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A3 (.DIODE(_2336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__B (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A1 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__B (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__B (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__B (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__B (.DIODE(_2351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A3 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A3 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A3 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A3 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A3 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A3 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A3 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A3 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A3 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A3 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__B (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__B (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__B (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__B (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__B (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__B (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__B (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__B (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__B (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__B (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__B (.DIODE(_2367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__B (.DIODE(_2367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A_N (.DIODE(_2367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__B (.DIODE(_2367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__B (.DIODE(_2367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A2 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A2 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A2 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__A2 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A2 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A2 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A2 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A2 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A2 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A2 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__C (.DIODE(_2373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__C (.DIODE(_2373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__C (.DIODE(_2373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__C (.DIODE(_2373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__C (.DIODE(_2373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__C (.DIODE(_2373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__C (.DIODE(_2373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__C (.DIODE(_2373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__C (.DIODE(_2373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__C (.DIODE(_2373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A (.DIODE(_2384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__B (.DIODE(_2388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__B (.DIODE(_2388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__B (.DIODE(_2388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__B (.DIODE(_2388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A2 (.DIODE(_2390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__A2 (.DIODE(_2390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A2 (.DIODE(_2390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A2 (.DIODE(_2390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A2 (.DIODE(_2390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A2 (.DIODE(_2390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A2 (.DIODE(_2390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A2 (.DIODE(_2390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A2 (.DIODE(_2390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A2 (.DIODE(_2390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__C (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__C (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__C (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__C (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__C (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__C (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__C (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__C (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__C (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__C (.DIODE(_2392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A (.DIODE(_2400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A (.DIODE(_2400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A (.DIODE(_2400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A (.DIODE(_2400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A (.DIODE(_2400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A (.DIODE(_2400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A (.DIODE(_2400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A (.DIODE(_2400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A (.DIODE(_2400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A (.DIODE(_2400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__B (.DIODE(_2407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__B (.DIODE(_2407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__B (.DIODE(_2407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__B (.DIODE(_2407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A2 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A2 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A2 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A2 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A2 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A2 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A2 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A2 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A2 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A2 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__C (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__C (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__C (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__C (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__C (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__C (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__C (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__C (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__C (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__C (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A2 (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A2 (.DIODE(_2433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__B1 (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__B1 (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__B (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__B (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__B (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__B (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__C (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__C (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__C (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__C (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__C (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__C (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__C (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__C (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__C (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__C (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__A (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A2 (.DIODE(_2462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__C (.DIODE(_2464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__C (.DIODE(_2464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__C (.DIODE(_2464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__C (.DIODE(_2464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__C (.DIODE(_2464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__C (.DIODE(_2464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__C (.DIODE(_2464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__C (.DIODE(_2464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__C (.DIODE(_2464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__C (.DIODE(_2464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__A (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__A (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A3 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A3 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A3 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A3 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A3 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A3 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A3 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A3 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A3 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A3 (.DIODE(_2480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__B (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__B (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__B (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__B (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__B (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__B (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__B (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__B (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__B (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__B (.DIODE(_2482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A1 (.DIODE(_2489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A1 (.DIODE(_2489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A1 (.DIODE(_2489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A1 (.DIODE(_2489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A1 (.DIODE(_2489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A1 (.DIODE(_2489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A1 (.DIODE(_2489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A1 (.DIODE(_2489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(_2489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A1 (.DIODE(_2489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A3 (.DIODE(_2495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A3 (.DIODE(_2495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A3 (.DIODE(_2495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A3 (.DIODE(_2495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A3 (.DIODE(_2495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A3 (.DIODE(_2495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A3 (.DIODE(_2495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A3 (.DIODE(_2495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A3 (.DIODE(_2495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A3 (.DIODE(_2495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__B (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__B (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__B (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__B (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__B (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__B (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__B (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__B (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__B (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__B (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A1 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A1 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A1 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A1 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A1 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A1 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A1 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A1 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A1 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A1 (.DIODE(_2503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A3 (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A3 (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A3 (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A3 (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A3 (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A3 (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A3 (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A3 (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A3 (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A3 (.DIODE(_2510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__B (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__B (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__B (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__B (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__B (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__B (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__B (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__B (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__B (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A1 (.DIODE(_2517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A1 (.DIODE(_2517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A1 (.DIODE(_2517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A1 (.DIODE(_2517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A1 (.DIODE(_2517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A1 (.DIODE(_2517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A1 (.DIODE(_2517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A1 (.DIODE(_2517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A1 (.DIODE(_2517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A1 (.DIODE(_2517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A3 (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A3 (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A3 (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A3 (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A3 (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A3 (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A3 (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A3 (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A3 (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A3 (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__B (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__B (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__B (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__B (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__B (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__B (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__B (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__B (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__B (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__B (.DIODE(_2527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A1 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A1 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A1 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A1 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A1 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A1 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A1 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A1 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A1 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A1 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__B (.DIODE(_2539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__B (.DIODE(_2539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__B (.DIODE(_2539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__B (.DIODE(_2539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A3 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A3 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A3 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A3 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A3 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A3 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A3 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A3 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A3 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A3 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B (.DIODE(_2543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__B (.DIODE(_2543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__B (.DIODE(_2543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__B (.DIODE(_2543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__B (.DIODE(_2543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__B (.DIODE(_2543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__B (.DIODE(_2543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__B (.DIODE(_2543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__B (.DIODE(_2543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__B (.DIODE(_2543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A1 (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A1 (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A1 (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A1 (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A1 (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A1 (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A1 (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A1 (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A1 (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A1 (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__B (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__B (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__B (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__B (.DIODE(_2555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A3 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A3 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A3 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A3 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A3 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A3 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A3 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A3 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A3 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A3 (.DIODE(_2557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__B (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__B (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__B (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__B (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__B (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__B (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__B (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__B (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__B (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__B (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__B (.DIODE(_2572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__B (.DIODE(_2572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__B (.DIODE(_2572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__B (.DIODE(_2572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A3 (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A3 (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A3 (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A3 (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A3 (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A3 (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A3 (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A3 (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A3 (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A3 (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__A1 (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A1 (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A1 (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A1 (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A1 (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A1 (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A1 (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A1 (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A1 (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A1 (.DIODE(_2576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A1 (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A1 (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A1 (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A1 (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A1 (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A1 (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A1 (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A1 (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A1 (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A1 (.DIODE(_2588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__B (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__B (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__B (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__B (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A3 (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A3 (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A3 (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A3 (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A3 (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A3 (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A3 (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A3 (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A3 (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A3 (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__B (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__B (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__B (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__B (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__B (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__B (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__B (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__B (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__B (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__B (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A1 (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__B (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__B (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__B (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__B (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A3 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A3 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A3 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A3 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A3 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A3 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A3 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A3 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A3 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A3 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__A1 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A1 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A1 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A1 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A1 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A1 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A1 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A1 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A1 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A1 (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__B (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__B (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__B (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A2 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A2 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A2 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A2 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A2 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A2 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A2 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A2 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A2 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A2 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__B1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__B1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__B1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__B1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__B1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__B1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__B1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__B1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__B1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B1 (.DIODE(_2625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A2 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A2 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A2 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A2 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A2 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A2 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A2 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A2 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A2 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A2 (.DIODE(_2632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__C (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__C (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__C (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__C (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__C (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__C (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__C (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__C (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__C (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__C (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__A (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A2 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A2 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A2 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A2 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A2 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A2 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A2 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A2 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A2 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A2 (.DIODE(_2650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__C (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__C (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__C (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__C (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__C (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__C (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__C (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__C (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__C (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__C (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__C (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__C (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__C (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__C (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__C (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__C (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__C (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__C (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__C (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__C (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__C (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__C (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__C (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__A (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A (.DIODE(_2681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__S (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__S (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__S (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__S (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__S (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__S (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__S (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__S (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__C (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__C (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__C (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__C (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__C (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__C (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__C (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__C (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__C (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__C (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__A (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__A (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__S (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__S (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__S (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__S (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__S (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__S (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__S (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__S (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A2 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A2 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A2 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__A2 (.DIODE(_2730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A2 (.DIODE(_2730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A2 (.DIODE(_2730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A2 (.DIODE(_2730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A2 (.DIODE(_2730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A2 (.DIODE(_2730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A2 (.DIODE(_2730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A2 (.DIODE(_2730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A2 (.DIODE(_2730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A2 (.DIODE(_2730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__C (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__C (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__C (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__A (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__C (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__C (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__C (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__C (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__C (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__C (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__C (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__C (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__C (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__C (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A2 (.DIODE(_2747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A2 (.DIODE(_2747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A2 (.DIODE(_2747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A (.DIODE(_2747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A2 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A2 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A2 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A2 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A2 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A2 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A2 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A2 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A2 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A2 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__A (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__A (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__C (.DIODE(_2750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__C (.DIODE(_2750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__C (.DIODE(_2750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A (.DIODE(_2750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__C (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__C (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__C (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__C (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__C (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__C (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__C (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__C (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__C (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__C (.DIODE(_2751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__A (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A (.DIODE(_2762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__A (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__A (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__A (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__A (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__A (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A3 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A3 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__A3 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A3 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A3 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A3 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A3 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A3 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A3 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A3 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__B (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A (.DIODE(_2791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__A (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__A (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__A (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__A (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__A (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__A (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__A (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__A (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A (.DIODE(_2793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__A (.DIODE(_2795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__A (.DIODE(_2795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A (.DIODE(_2795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A (.DIODE(_2795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__A (.DIODE(_2795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A (.DIODE(_2795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A (.DIODE(_2795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__A (.DIODE(_2795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A (.DIODE(_2795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A (.DIODE(_2795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__A (.DIODE(_2797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__A (.DIODE(_2797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A (.DIODE(_2797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__A (.DIODE(_2797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A (.DIODE(_2797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A (.DIODE(_2797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A (.DIODE(_2797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__A (.DIODE(_2797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A (.DIODE(_2797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A (.DIODE(_2797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__A (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__A (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__A (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__A (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__A (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__A (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__A (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__A (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__A (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__A (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__A (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A (.DIODE(_2803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__C (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__C (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__C (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__C (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__C (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__C (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__C (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__C (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__C (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__C (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A2 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A2 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A2 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__A2 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A2 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A2 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A2 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A2 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A2 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A2 (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__C (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__C (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__C (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__C (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__C (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__C (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__C (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__C (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__C (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__C (.DIODE(_2832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__A (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__A (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__A (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__A (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__A (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__S (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A3 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A3 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A3 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A3 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A3 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A3 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A3 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A3 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__A3 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A3 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__B (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__B (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__B (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__B (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__B (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__B (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__B (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__B (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__B (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__B (.DIODE(_2861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A1 (.DIODE(_2867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A3 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__A3 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__A3 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A3 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A3 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__A3 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__A3 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__A3 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__A3 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__A3 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A3 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A3 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A3 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__A (.DIODE(_2879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__B (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__B (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__B (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__A (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__B (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__B (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__B (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__B (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__B (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__B (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__B (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__B (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__B (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__B (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__A1 (.DIODE(_2884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__A1 (.DIODE(_2884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A1 (.DIODE(_2884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A1 (.DIODE(_2884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__A1 (.DIODE(_2884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__A1 (.DIODE(_2884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__A1 (.DIODE(_2884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__A1 (.DIODE(_2884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__A1 (.DIODE(_2884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A1 (.DIODE(_2884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__A (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__A (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__A (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__A (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__A (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__A (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A (.DIODE(_2895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__A (.DIODE(_2895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__A (.DIODE(_2895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A (.DIODE(_2895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__A (.DIODE(_2895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__A (.DIODE(_2895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__A (.DIODE(_2895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__A (.DIODE(_2895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__A (.DIODE(_2895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__A (.DIODE(_2895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__A1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__A1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A1 (.DIODE(_2898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A3 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A3 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A3 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A3 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A3 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A3 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__A3 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__A3 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A3 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A3 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__B (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__B (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__B (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__B (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__B (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__B (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__B (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__B (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__B (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__B (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__A (.DIODE(_2919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__A (.DIODE(_2919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__A (.DIODE(_2919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__A (.DIODE(_2919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__A (.DIODE(_2919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__A (.DIODE(_2919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__A (.DIODE(_2919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__A (.DIODE(_2919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__A (.DIODE(_2919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__A (.DIODE(_2919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A3 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A3 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A3 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__A3 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__A3 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__A3 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__A3 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A3 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__A3 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A3 (.DIODE(_2922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__B (.DIODE(_2924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__B (.DIODE(_2924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__B (.DIODE(_2924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__B (.DIODE(_2924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__B (.DIODE(_2924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__B (.DIODE(_2924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__B (.DIODE(_2924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__B (.DIODE(_2924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__B (.DIODE(_2924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__B (.DIODE(_2924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6280__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__A (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__A1 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A1 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__A1 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A1 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A1 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A1 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A1 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A1 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A1 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__A1 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__A3 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A3 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A3 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A3 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__A3 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__A3 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A3 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__A3 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A3 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__A3 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__B (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__B (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__B (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__B (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__B (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__B (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__B (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__B (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__B (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__B (.DIODE(_2944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A2 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A2 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__A2 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A2 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A2 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A2 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__A2 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__A2 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A2 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A2 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__C (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__C (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__C (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__C (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__C (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__C (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__C (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__C (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__C (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__C (.DIODE(_2962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__A (.DIODE(_2971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__A (.DIODE(_2971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__A (.DIODE(_2971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__A (.DIODE(_2971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__A (.DIODE(_2971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__A (.DIODE(_2971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A (.DIODE(_2971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__A (.DIODE(_2971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__A (.DIODE(_2971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__A (.DIODE(_2971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A1 (.DIODE(_2977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A1 (.DIODE(_2977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A1 (.DIODE(_2977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A1 (.DIODE(_2977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A1 (.DIODE(_2977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__A1 (.DIODE(_2977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A1 (.DIODE(_2977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A1 (.DIODE(_2977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__A1 (.DIODE(_2977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A1 (.DIODE(_2977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A3 (.DIODE(_2980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__A3 (.DIODE(_2980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__A3 (.DIODE(_2980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A (.DIODE(_2980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A3 (.DIODE(_2981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A3 (.DIODE(_2981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A3 (.DIODE(_2981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A3 (.DIODE(_2981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A3 (.DIODE(_2981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__A3 (.DIODE(_2981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A3 (.DIODE(_2981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A3 (.DIODE(_2981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__A3 (.DIODE(_2981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A3 (.DIODE(_2981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__B (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__B (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__B (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__B (.DIODE(_2983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__B (.DIODE(_2983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__B (.DIODE(_2983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__B (.DIODE(_2983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__B (.DIODE(_2983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__B (.DIODE(_2983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__B (.DIODE(_2983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__B (.DIODE(_2983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__B (.DIODE(_2983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__B (.DIODE(_2983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__A1 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A1 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__A1 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__A1 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__A1 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__A1 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A1 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A1 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__A1 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__A1 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A3 (.DIODE(_3000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__A3 (.DIODE(_3000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A3 (.DIODE(_3000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__A3 (.DIODE(_3000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A3 (.DIODE(_3000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__A3 (.DIODE(_3000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__A3 (.DIODE(_3000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__A3 (.DIODE(_3000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__A3 (.DIODE(_3000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A3 (.DIODE(_3000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A1 (.DIODE(_3010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A3 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__A3 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__A3 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__A (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A3 (.DIODE(_3019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A3 (.DIODE(_3019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A3 (.DIODE(_3019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__A3 (.DIODE(_3019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6237__A3 (.DIODE(_3019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A3 (.DIODE(_3019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A3 (.DIODE(_3019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A3 (.DIODE(_3019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__A3 (.DIODE(_3019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A3 (.DIODE(_3019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__B (.DIODE(_3020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__B (.DIODE(_3020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__B (.DIODE(_3020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A (.DIODE(_3020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__B (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__B (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__B (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__B (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__B (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__B (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__B (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__B (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__B (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__B (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6258__A1 (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A1 (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__A1 (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__A1 (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A1 (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A1 (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A1 (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__A1 (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6237__A1 (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A1 (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A3 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A3 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__A3 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A3 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__A3 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__A3 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__A3 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A3 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__A3 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6258__A3 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__B (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__B (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__B (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__B (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__B (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__B (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__B (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__B (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__B (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__B (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__A1 (.DIODE(_3042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A1 (.DIODE(_3042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A1 (.DIODE(_3042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__A1 (.DIODE(_3042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A1 (.DIODE(_3042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__A1 (.DIODE(_3042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__A1 (.DIODE(_3042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__A1 (.DIODE(_3042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A1 (.DIODE(_3042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__A1 (.DIODE(_3042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__A3 (.DIODE(_3057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__A3 (.DIODE(_3057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A3 (.DIODE(_3057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__A (.DIODE(_3057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A3 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__A3 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A3 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A3 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A3 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A3 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A3 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__A3 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A3 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__A3 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__B (.DIODE(_3059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__B (.DIODE(_3059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__B (.DIODE(_3059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__A (.DIODE(_3059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__B (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__B (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__B (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__B (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__B (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__B (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__B (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__B (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__B (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__B (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__A1 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A1 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A1 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__A1 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A1 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__A1 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__A1 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A1 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A1 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__A1 (.DIODE(_3069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__A3 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__A3 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A3 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A3 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__A3 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__A3 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A3 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A3 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__A3 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A3 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__B (.DIODE(_3079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__A1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A3 (.DIODE(_3096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A3 (.DIODE(_3096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A3 (.DIODE(_3096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A3 (.DIODE(_3096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A3 (.DIODE(_3096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A3 (.DIODE(_3096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A3 (.DIODE(_3096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A3 (.DIODE(_3096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A3 (.DIODE(_3096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__A3 (.DIODE(_3096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__B (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__B (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__B (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__B (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__B (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__B (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__B (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__B (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__B (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__B (.DIODE(_3098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6378__A1 (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A1 (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A1 (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A1 (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A1 (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A1 (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A1 (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A1 (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A1 (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A1 (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__A1 (.DIODE(_3112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__A1 (.DIODE(_3112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A1 (.DIODE(_3112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__A1 (.DIODE(_3112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A1 (.DIODE(_3112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__A1 (.DIODE(_3112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A1 (.DIODE(_3112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A1 (.DIODE(_3112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__A1 (.DIODE(_3112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A1 (.DIODE(_3112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A3 (.DIODE(_3115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A3 (.DIODE(_3115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A3 (.DIODE(_3115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A (.DIODE(_3115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__A3 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__A3 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__A3 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A3 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__A3 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A3 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__A3 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A3 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A3 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__A3 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__B (.DIODE(_3117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__B (.DIODE(_3117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__B (.DIODE(_3117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__A (.DIODE(_3117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__B (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__B (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__B (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__B (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__B (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__B (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__B (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__B (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__B (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__B (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__A1 (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A1 (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__A1 (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A1 (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__A1 (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A1 (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A1 (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A1 (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A1 (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__A1 (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A3 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A3 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__A3 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__A3 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__A3 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A3 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A3 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__A3 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A3 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__A3 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A3 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__A3 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A3 (.DIODE(_3135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__B (.DIODE(_3136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__B (.DIODE(_3136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__B (.DIODE(_3136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A (.DIODE(_3136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__B (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__B (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__B (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__B (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__B (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__B (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__B (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__B (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__B (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__B (.DIODE(_3137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__A2 (.DIODE(_3157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A2 (.DIODE(_3157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__A2 (.DIODE(_3157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A2 (.DIODE(_3157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__A2 (.DIODE(_3157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__A2 (.DIODE(_3157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A2 (.DIODE(_3157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A2 (.DIODE(_3157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__A2 (.DIODE(_3157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__A2 (.DIODE(_3157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__C (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__C (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__C (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__C (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__C (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__C (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__C (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__C (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__C (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__C (.DIODE(_3159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__S (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__S (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__S (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__S (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__S (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__S (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__S (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__S (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(c0_o_c_data_page));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(c0_o_c_instr_long));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(c0_o_c_instr_page));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(c0_o_icache_flush));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(c0_o_instr_long_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(c0_o_instr_long_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(c0_o_instr_long_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(c0_o_instr_long_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(c0_o_instr_long_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(c0_o_instr_long_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(c0_o_instr_long_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(c0_o_instr_long_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(c0_o_mem_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(c0_o_mem_addr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(c0_o_mem_addr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(c0_o_mem_addr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(c0_o_mem_addr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(c0_o_mem_addr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(c0_o_mem_addr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(c0_o_mem_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(c0_o_mem_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(c0_o_mem_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(c0_o_mem_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(c0_o_mem_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(c0_o_mem_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(c0_o_mem_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(c0_o_mem_addr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(c0_o_mem_addr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(c0_o_mem_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(c0_o_mem_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(c0_o_mem_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(c0_o_mem_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(c0_o_mem_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(c0_o_mem_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(c0_o_mem_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(c0_o_mem_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(c0_o_mem_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(c0_o_mem_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(c0_o_mem_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(c0_o_mem_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(c0_o_mem_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(c0_o_mem_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(c0_o_mem_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(c0_o_mem_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(c0_o_mem_high_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(c0_o_mem_high_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(c0_o_mem_high_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(c0_o_mem_high_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(c0_o_mem_high_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(c0_o_mem_high_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(c0_o_mem_high_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(c0_o_mem_high_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(c0_o_mem_long_mode));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(c0_o_mem_req));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(c0_o_mem_sel[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(c0_o_mem_sel[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(c0_o_mem_we));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(c0_o_req_active));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(c0_o_req_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(c0_o_req_addr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(c0_o_req_addr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(c0_o_req_addr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(c0_o_req_addr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(c0_o_req_addr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(c0_o_req_addr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(c0_o_req_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(c0_o_req_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(c0_o_req_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(c0_o_req_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(c0_o_req_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(c0_o_req_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(c0_o_req_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(c0_o_req_addr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(c0_o_req_addr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(c0_o_req_ppl_submit));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(c0_sr_bus_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(c0_sr_bus_addr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(c0_sr_bus_addr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(c0_sr_bus_addr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(c0_sr_bus_addr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(c0_sr_bus_addr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(c0_sr_bus_addr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(c0_sr_bus_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(c0_sr_bus_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(c0_sr_bus_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(c0_sr_bus_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(c0_sr_bus_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(c0_sr_bus_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(c0_sr_bus_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(c0_sr_bus_addr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(c0_sr_bus_addr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(c0_sr_bus_data_o[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(c0_sr_bus_data_o[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(c0_sr_bus_data_o[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(c0_sr_bus_data_o[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(c0_sr_bus_data_o[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(c0_sr_bus_data_o[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(c0_sr_bus_data_o[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(c0_sr_bus_data_o[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(c0_sr_bus_data_o[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input101_A (.DIODE(c0_sr_bus_data_o[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input102_A (.DIODE(c0_sr_bus_data_o[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input103_A (.DIODE(c0_sr_bus_data_o[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input104_A (.DIODE(c0_sr_bus_data_o[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input105_A (.DIODE(c0_sr_bus_we));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__CLK (.DIODE(clknet_leaf_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__CLK (.DIODE(clknet_leaf_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__CLK (.DIODE(clknet_leaf_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__CLK (.DIODE(clknet_leaf_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__CLK (.DIODE(clknet_leaf_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__CLK (.DIODE(clknet_leaf_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__CLK (.DIODE(clknet_leaf_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__CLK (.DIODE(clknet_leaf_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__CLK (.DIODE(clknet_leaf_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_input106_A (.DIODE(c1_o_c_data_page));
 sky130_fd_sc_hd__diode_2 ANTENNA_input107_A (.DIODE(c1_o_c_instr_long));
 sky130_fd_sc_hd__diode_2 ANTENNA_input108_A (.DIODE(c1_o_c_instr_page));
 sky130_fd_sc_hd__diode_2 ANTENNA_input109_A (.DIODE(c1_o_icache_flush));
 sky130_fd_sc_hd__diode_2 ANTENNA_input110_A (.DIODE(c1_o_instr_long_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input111_A (.DIODE(c1_o_instr_long_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input112_A (.DIODE(c1_o_instr_long_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input113_A (.DIODE(c1_o_instr_long_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input114_A (.DIODE(c1_o_instr_long_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input115_A (.DIODE(c1_o_instr_long_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input116_A (.DIODE(c1_o_instr_long_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input117_A (.DIODE(c1_o_instr_long_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input118_A (.DIODE(c1_o_mem_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input119_A (.DIODE(c1_o_mem_addr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input120_A (.DIODE(c1_o_mem_addr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input121_A (.DIODE(c1_o_mem_addr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input122_A (.DIODE(c1_o_mem_addr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input123_A (.DIODE(c1_o_mem_addr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input124_A (.DIODE(c1_o_mem_addr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input125_A (.DIODE(c1_o_mem_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input126_A (.DIODE(c1_o_mem_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input127_A (.DIODE(c1_o_mem_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input128_A (.DIODE(c1_o_mem_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input129_A (.DIODE(c1_o_mem_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input130_A (.DIODE(c1_o_mem_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input131_A (.DIODE(c1_o_mem_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input132_A (.DIODE(c1_o_mem_addr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input133_A (.DIODE(c1_o_mem_addr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input134_A (.DIODE(c1_o_mem_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input135_A (.DIODE(c1_o_mem_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input136_A (.DIODE(c1_o_mem_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input137_A (.DIODE(c1_o_mem_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input138_A (.DIODE(c1_o_mem_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input139_A (.DIODE(c1_o_mem_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input140_A (.DIODE(c1_o_mem_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input141_A (.DIODE(c1_o_mem_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input142_A (.DIODE(c1_o_mem_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input143_A (.DIODE(c1_o_mem_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input144_A (.DIODE(c1_o_mem_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input145_A (.DIODE(c1_o_mem_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input146_A (.DIODE(c1_o_mem_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input147_A (.DIODE(c1_o_mem_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input148_A (.DIODE(c1_o_mem_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input149_A (.DIODE(c1_o_mem_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input150_A (.DIODE(c1_o_mem_high_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input151_A (.DIODE(c1_o_mem_high_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input152_A (.DIODE(c1_o_mem_high_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input153_A (.DIODE(c1_o_mem_high_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input154_A (.DIODE(c1_o_mem_high_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input155_A (.DIODE(c1_o_mem_high_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input156_A (.DIODE(c1_o_mem_high_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input157_A (.DIODE(c1_o_mem_high_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input158_A (.DIODE(c1_o_mem_long_mode));
 sky130_fd_sc_hd__diode_2 ANTENNA_input159_A (.DIODE(c1_o_mem_req));
 sky130_fd_sc_hd__diode_2 ANTENNA_input160_A (.DIODE(c1_o_mem_sel[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input161_A (.DIODE(c1_o_mem_sel[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input162_A (.DIODE(c1_o_mem_we));
 sky130_fd_sc_hd__diode_2 ANTENNA_input163_A (.DIODE(c1_o_req_active));
 sky130_fd_sc_hd__diode_2 ANTENNA_input164_A (.DIODE(c1_o_req_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input165_A (.DIODE(c1_o_req_addr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input166_A (.DIODE(c1_o_req_addr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input167_A (.DIODE(c1_o_req_addr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input168_A (.DIODE(c1_o_req_addr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input169_A (.DIODE(c1_o_req_addr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input170_A (.DIODE(c1_o_req_addr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input171_A (.DIODE(c1_o_req_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input172_A (.DIODE(c1_o_req_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input173_A (.DIODE(c1_o_req_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input174_A (.DIODE(c1_o_req_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input175_A (.DIODE(c1_o_req_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input176_A (.DIODE(c1_o_req_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input177_A (.DIODE(c1_o_req_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input178_A (.DIODE(c1_o_req_addr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input179_A (.DIODE(c1_o_req_addr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input180_A (.DIODE(c1_o_req_ppl_submit));
 sky130_fd_sc_hd__diode_2 ANTENNA_input181_A (.DIODE(c1_sr_bus_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input182_A (.DIODE(c1_sr_bus_addr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input183_A (.DIODE(c1_sr_bus_addr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input184_A (.DIODE(c1_sr_bus_addr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input185_A (.DIODE(c1_sr_bus_addr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input186_A (.DIODE(c1_sr_bus_addr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input187_A (.DIODE(c1_sr_bus_addr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input188_A (.DIODE(c1_sr_bus_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input189_A (.DIODE(c1_sr_bus_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input190_A (.DIODE(c1_sr_bus_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input191_A (.DIODE(c1_sr_bus_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input192_A (.DIODE(c1_sr_bus_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input193_A (.DIODE(c1_sr_bus_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input194_A (.DIODE(c1_sr_bus_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input195_A (.DIODE(c1_sr_bus_addr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input196_A (.DIODE(c1_sr_bus_addr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input197_A (.DIODE(c1_sr_bus_data_o[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input198_A (.DIODE(c1_sr_bus_data_o[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input199_A (.DIODE(c1_sr_bus_data_o[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input200_A (.DIODE(c1_sr_bus_data_o[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input201_A (.DIODE(c1_sr_bus_data_o[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input202_A (.DIODE(c1_sr_bus_data_o[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input203_A (.DIODE(c1_sr_bus_data_o[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input204_A (.DIODE(c1_sr_bus_data_o[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input205_A (.DIODE(c1_sr_bus_data_o[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input206_A (.DIODE(c1_sr_bus_data_o[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input207_A (.DIODE(c1_sr_bus_data_o[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input208_A (.DIODE(c1_sr_bus_data_o[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input209_A (.DIODE(c1_sr_bus_data_o[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input210_A (.DIODE(c1_sr_bus_we));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_core_clock_A (.DIODE(core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_input211_A (.DIODE(core_reset));
 sky130_fd_sc_hd__diode_2 ANTENNA_input212_A (.DIODE(dcache_mem_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA_input213_A (.DIODE(dcache_mem_exception));
 sky130_fd_sc_hd__diode_2 ANTENNA_input214_A (.DIODE(dcache_mem_o_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input215_A (.DIODE(dcache_mem_o_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input216_A (.DIODE(dcache_mem_o_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input217_A (.DIODE(dcache_mem_o_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input218_A (.DIODE(dcache_mem_o_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input219_A (.DIODE(dcache_mem_o_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input220_A (.DIODE(dcache_mem_o_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input221_A (.DIODE(dcache_mem_o_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input222_A (.DIODE(dcache_mem_o_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input223_A (.DIODE(dcache_mem_o_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input224_A (.DIODE(dcache_mem_o_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input225_A (.DIODE(dcache_mem_o_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input226_A (.DIODE(dcache_mem_o_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input227_A (.DIODE(dcache_mem_o_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input228_A (.DIODE(dcache_mem_o_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input229_A (.DIODE(dcache_mem_o_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input230_A (.DIODE(dcache_wb_4_burst));
 sky130_fd_sc_hd__diode_2 ANTENNA_input231_A (.DIODE(dcache_wb_adr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input232_A (.DIODE(dcache_wb_adr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input233_A (.DIODE(dcache_wb_adr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input234_A (.DIODE(dcache_wb_adr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input235_A (.DIODE(dcache_wb_adr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input236_A (.DIODE(dcache_wb_adr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input237_A (.DIODE(dcache_wb_adr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input238_A (.DIODE(dcache_wb_adr[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input239_A (.DIODE(dcache_wb_adr[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input240_A (.DIODE(dcache_wb_adr[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input241_A (.DIODE(dcache_wb_adr[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input242_A (.DIODE(dcache_wb_adr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input243_A (.DIODE(dcache_wb_adr[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input244_A (.DIODE(dcache_wb_adr[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input245_A (.DIODE(dcache_wb_adr[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input246_A (.DIODE(dcache_wb_adr[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input247_A (.DIODE(dcache_wb_adr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input248_A (.DIODE(dcache_wb_adr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input249_A (.DIODE(dcache_wb_adr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input250_A (.DIODE(dcache_wb_adr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input251_A (.DIODE(dcache_wb_adr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input252_A (.DIODE(dcache_wb_adr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input253_A (.DIODE(dcache_wb_adr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input254_A (.DIODE(dcache_wb_adr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input255_A (.DIODE(dcache_wb_cyc));
 sky130_fd_sc_hd__diode_2 ANTENNA_input256_A (.DIODE(dcache_wb_o_dat[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input257_A (.DIODE(dcache_wb_o_dat[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input258_A (.DIODE(dcache_wb_o_dat[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input259_A (.DIODE(dcache_wb_o_dat[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input260_A (.DIODE(dcache_wb_o_dat[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input261_A (.DIODE(dcache_wb_o_dat[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input262_A (.DIODE(dcache_wb_o_dat[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input263_A (.DIODE(dcache_wb_o_dat[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input264_A (.DIODE(dcache_wb_o_dat[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input265_A (.DIODE(dcache_wb_o_dat[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input266_A (.DIODE(dcache_wb_o_dat[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input267_A (.DIODE(dcache_wb_o_dat[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input268_A (.DIODE(dcache_wb_o_dat[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input269_A (.DIODE(dcache_wb_o_dat[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input270_A (.DIODE(dcache_wb_o_dat[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input271_A (.DIODE(dcache_wb_o_dat[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input272_A (.DIODE(dcache_wb_sel[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input273_A (.DIODE(dcache_wb_sel[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input274_A (.DIODE(dcache_wb_stb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input275_A (.DIODE(dcache_wb_we));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__B (.DIODE(\dmmu0.page_table[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__A1 (.DIODE(\dmmu0.page_table[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__B (.DIODE(\dmmu0.page_table[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__A1 (.DIODE(\dmmu0.page_table[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__B (.DIODE(\dmmu0.page_table[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__A1 (.DIODE(\dmmu0.page_table[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__B (.DIODE(\dmmu0.page_table[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A1 (.DIODE(\dmmu0.page_table[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__B (.DIODE(\dmmu0.page_table[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__A1 (.DIODE(\dmmu0.page_table[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__B (.DIODE(\dmmu0.page_table[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__A3 (.DIODE(\dmmu0.page_table[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__B (.DIODE(\dmmu0.page_table[3][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A1 (.DIODE(\dmmu0.page_table[3][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__B (.DIODE(\dmmu0.page_table[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__A1 (.DIODE(\dmmu0.page_table[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__B (.DIODE(\dmmu0.page_table[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__A3 (.DIODE(\dmmu0.page_table[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__B (.DIODE(\dmmu0.page_table[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A3 (.DIODE(\dmmu0.page_table[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__B (.DIODE(\dmmu0.page_table[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__A1 (.DIODE(\dmmu0.page_table[3][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__B (.DIODE(\dmmu0.page_table[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A1 (.DIODE(\dmmu0.page_table[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__B (.DIODE(\dmmu0.page_table[6][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A0 (.DIODE(\dmmu0.page_table[6][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__B (.DIODE(\dmmu0.page_table[9][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A1 (.DIODE(\dmmu0.page_table[9][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__B (.DIODE(\dmmu0.page_table[9][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__A1 (.DIODE(\dmmu0.page_table[9][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__B (.DIODE(\dmmu0.page_table[9][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A1 (.DIODE(\dmmu0.page_table[9][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input276_A (.DIODE(ic0_mem_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA_input277_A (.DIODE(ic0_mem_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input278_A (.DIODE(ic0_mem_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input279_A (.DIODE(ic0_mem_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input280_A (.DIODE(ic0_mem_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input281_A (.DIODE(ic0_mem_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input282_A (.DIODE(ic0_mem_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input283_A (.DIODE(ic0_mem_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input284_A (.DIODE(ic0_mem_data[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input285_A (.DIODE(ic0_mem_data[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input286_A (.DIODE(ic0_mem_data[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input287_A (.DIODE(ic0_mem_data[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input288_A (.DIODE(ic0_mem_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input289_A (.DIODE(ic0_mem_data[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input290_A (.DIODE(ic0_mem_data[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input291_A (.DIODE(ic0_mem_data[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input292_A (.DIODE(ic0_mem_data[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input293_A (.DIODE(ic0_mem_data[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input294_A (.DIODE(ic0_mem_data[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input295_A (.DIODE(ic0_mem_data[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input296_A (.DIODE(ic0_mem_data[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input297_A (.DIODE(ic0_mem_data[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input298_A (.DIODE(ic0_mem_data[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input299_A (.DIODE(ic0_mem_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input300_A (.DIODE(ic0_mem_data[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input301_A (.DIODE(ic0_mem_data[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input302_A (.DIODE(ic0_mem_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input303_A (.DIODE(ic0_mem_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input304_A (.DIODE(ic0_mem_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input305_A (.DIODE(ic0_mem_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input306_A (.DIODE(ic0_mem_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input307_A (.DIODE(ic0_mem_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input308_A (.DIODE(ic0_mem_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input309_A (.DIODE(ic0_wb_adr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input310_A (.DIODE(ic0_wb_adr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input311_A (.DIODE(ic0_wb_adr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input312_A (.DIODE(ic0_wb_adr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input313_A (.DIODE(ic0_wb_adr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input314_A (.DIODE(ic0_wb_adr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input315_A (.DIODE(ic0_wb_adr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input316_A (.DIODE(ic0_wb_adr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input317_A (.DIODE(ic0_wb_adr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input318_A (.DIODE(ic0_wb_adr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input319_A (.DIODE(ic0_wb_adr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input320_A (.DIODE(ic0_wb_adr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input321_A (.DIODE(ic0_wb_adr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input322_A (.DIODE(ic0_wb_adr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input323_A (.DIODE(ic0_wb_adr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input324_A (.DIODE(ic0_wb_adr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input325_A (.DIODE(ic0_wb_cyc));
 sky130_fd_sc_hd__diode_2 ANTENNA_input326_A (.DIODE(ic0_wb_sel[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input327_A (.DIODE(ic0_wb_sel[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input328_A (.DIODE(ic0_wb_stb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input329_A (.DIODE(ic0_wb_we));
 sky130_fd_sc_hd__diode_2 ANTENNA_input330_A (.DIODE(ic1_mem_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA_input331_A (.DIODE(ic1_mem_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input332_A (.DIODE(ic1_mem_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input333_A (.DIODE(ic1_mem_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input334_A (.DIODE(ic1_mem_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input335_A (.DIODE(ic1_mem_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input336_A (.DIODE(ic1_mem_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input337_A (.DIODE(ic1_mem_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input338_A (.DIODE(ic1_mem_data[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input339_A (.DIODE(ic1_mem_data[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input340_A (.DIODE(ic1_mem_data[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input341_A (.DIODE(ic1_mem_data[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input342_A (.DIODE(ic1_mem_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input343_A (.DIODE(ic1_mem_data[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input344_A (.DIODE(ic1_mem_data[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input345_A (.DIODE(ic1_mem_data[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input346_A (.DIODE(ic1_mem_data[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input347_A (.DIODE(ic1_mem_data[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input348_A (.DIODE(ic1_mem_data[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input349_A (.DIODE(ic1_mem_data[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input350_A (.DIODE(ic1_mem_data[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input351_A (.DIODE(ic1_mem_data[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input352_A (.DIODE(ic1_mem_data[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input353_A (.DIODE(ic1_mem_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input354_A (.DIODE(ic1_mem_data[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input355_A (.DIODE(ic1_mem_data[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input356_A (.DIODE(ic1_mem_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input357_A (.DIODE(ic1_mem_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input358_A (.DIODE(ic1_mem_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input359_A (.DIODE(ic1_mem_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input360_A (.DIODE(ic1_mem_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input361_A (.DIODE(ic1_mem_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input362_A (.DIODE(ic1_mem_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input363_A (.DIODE(ic1_wb_adr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input364_A (.DIODE(ic1_wb_adr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input365_A (.DIODE(ic1_wb_adr[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input366_A (.DIODE(ic1_wb_adr[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input367_A (.DIODE(ic1_wb_adr[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input368_A (.DIODE(ic1_wb_adr[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input369_A (.DIODE(ic1_wb_adr[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input370_A (.DIODE(ic1_wb_adr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input371_A (.DIODE(ic1_wb_adr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input372_A (.DIODE(ic1_wb_adr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input373_A (.DIODE(ic1_wb_adr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input374_A (.DIODE(ic1_wb_adr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input375_A (.DIODE(ic1_wb_adr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input376_A (.DIODE(ic1_wb_adr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input377_A (.DIODE(ic1_wb_adr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input378_A (.DIODE(ic1_wb_adr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input379_A (.DIODE(ic1_wb_cyc));
 sky130_fd_sc_hd__diode_2 ANTENNA_input380_A (.DIODE(ic1_wb_sel[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input381_A (.DIODE(ic1_wb_sel[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input382_A (.DIODE(ic1_wb_stb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input383_A (.DIODE(ic1_wb_we));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A2 (.DIODE(\immu_0.page_table[15][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A3 (.DIODE(\immu_0.page_table[15][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A2 (.DIODE(\immu_0.page_table[8][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A2 (.DIODE(\immu_0.page_table[8][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A2 (.DIODE(\immu_0.page_table[8][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A0 (.DIODE(\immu_0.page_table[8][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A2 (.DIODE(\immu_0.page_table[8][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__A0 (.DIODE(\immu_0.page_table[8][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A2 (.DIODE(\immu_0.page_table[9][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A3 (.DIODE(\immu_0.page_table[9][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A2 (.DIODE(\immu_0.page_table[9][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__A1 (.DIODE(\immu_0.page_table[9][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A0 (.DIODE(\immu_1.high_addr_off[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__B (.DIODE(\immu_1.high_addr_off[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__B (.DIODE(\immu_1.high_addr_off[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__B2 (.DIODE(\immu_1.page_table[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A0 (.DIODE(\immu_1.page_table[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__B2 (.DIODE(\immu_1.page_table[0][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__A0 (.DIODE(\immu_1.page_table[0][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__B (.DIODE(\immu_1.page_table[14][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__A0 (.DIODE(\immu_1.page_table[14][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__B (.DIODE(\immu_1.page_table[7][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__A3 (.DIODE(\immu_1.page_table[7][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__B (.DIODE(\immu_1.page_table[9][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__A1 (.DIODE(\immu_1.page_table[9][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input384_A (.DIODE(inner_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA_input385_A (.DIODE(inner_embed_mode));
 sky130_fd_sc_hd__diode_2 ANTENNA_input386_A (.DIODE(inner_ext_irq));
 sky130_fd_sc_hd__diode_2 ANTENNA_input387_A (.DIODE(inner_wb_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A1 (.DIODE(\inner_wb_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__B1 (.DIODE(\inner_wb_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__A (.DIODE(\inner_wb_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__B1 (.DIODE(\inner_wb_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__A (.DIODE(\inner_wb_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__A (.DIODE(\inner_wb_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__A (.DIODE(\inner_wb_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A (.DIODE(\inner_wb_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__A (.DIODE(\inner_wb_arbiter.o_sel_sig ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input388_A (.DIODE(inner_wb_err));
 sky130_fd_sc_hd__diode_2 ANTENNA_input389_A (.DIODE(inner_wb_i_dat[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input390_A (.DIODE(inner_wb_i_dat[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input391_A (.DIODE(inner_wb_i_dat[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input392_A (.DIODE(inner_wb_i_dat[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input393_A (.DIODE(inner_wb_i_dat[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input394_A (.DIODE(inner_wb_i_dat[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input395_A (.DIODE(inner_wb_i_dat[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input396_A (.DIODE(inner_wb_i_dat[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input397_A (.DIODE(inner_wb_i_dat[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input398_A (.DIODE(inner_wb_i_dat[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input399_A (.DIODE(inner_wb_i_dat[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input400_A (.DIODE(inner_wb_i_dat[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input401_A (.DIODE(inner_wb_i_dat[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input402_A (.DIODE(inner_wb_i_dat[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input403_A (.DIODE(inner_wb_i_dat[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input404_A (.DIODE(inner_wb_i_dat[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__B1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__7452__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__S (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__S (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__S0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__S0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__S (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__S1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__S1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__S1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__S1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__S1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3308__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__C1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__C1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__3333__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__A_N (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7454__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7436__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7446__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__7447__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__7448__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__7449__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__7450__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7451__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7437__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__7438__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__7439__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__7440__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__7441__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__7442__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7443__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7444__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7445__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7453__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__D_N (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__C_N (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__7489__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__A0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__S0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__S0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__S0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__S1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__S1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__S1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__S1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3261__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__C1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__C1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__C1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__A0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__A0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__A0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__A0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__A0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__A0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__A0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A0 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__A0 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__D (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__C (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__D (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__C (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A0 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A0 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7491__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7473__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__7474__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__7490__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__B_N (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__B_N (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__D (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__B_N (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__C (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__B_N (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__B2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6281__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__B2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__D_N (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout710_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__7492__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__7416__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__B (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A0 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A0 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A0 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A0 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A0 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__B2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A2 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__B2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A0 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A0 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__A0 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A0 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A0 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__A0 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__B (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A0 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A0 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A0 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A0 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__A0 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A0 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A0 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__S (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__S (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__S (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__S (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__S (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__S (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__S0 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__S1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__S1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__S1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__B1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__C1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__B1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__S1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__B1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A0 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A0 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A0 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A0 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__A0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A0 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__B1_N (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__A0 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__A0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__A0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A0 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A0 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__7393__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__7394__A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__7395__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__7396__A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__7397__A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__7398__A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__7399__A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__7400__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__7401__A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__7402__A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__7403__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__7404__A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__7405__A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__7406__A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__7407__A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__7408__A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__7409__A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__7410__A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__7411__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__7412__A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__7385__A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__7413__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__7414__A (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__7386__A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__7387__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__7388__A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__7389__A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__7390__A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__7391__A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__7392__A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__S (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__S (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__S1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__C1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__B (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__B (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__C1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__A1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__S1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__C1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A1 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__A1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A1 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__7342__A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__B (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__A_N (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__B (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__C (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__C (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__B (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__C (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__C (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__7493__A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__7456__A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__7419__A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__7503__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__7466__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__7429__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__7504__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__7467__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__7430__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__7505__A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__7468__A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__7431__A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__7506__A (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__7469__A (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__7432__A (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__7507__A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__7470__A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__7433__A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__7508__A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__7471__A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__7434__A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__7494__A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__7457__A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__7420__A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__7495__A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__7458__A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__7421__A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__7496__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__7459__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__7422__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__7497__A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__7460__A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__7423__A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__7498__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__7461__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__7424__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__7499__A (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__7462__A (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__7425__A (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__7500__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__7463__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__7426__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__7501__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__7464__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__7427__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__7502__A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__7465__A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__7428__A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_output407_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7380__A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__7344__A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__B1_N (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_output408_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__7382__A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__7381__A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__B1_N (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_output409_A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_output429_A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_output430_A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_output431_A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_output432_A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_output433_A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_output434_A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_output435_A (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_output436_A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_output437_A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_output438_A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_output439_A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_output440_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_output441_A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_output442_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_output443_A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_output444_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_output445_A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_output446_A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_output447_A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_output448_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_output449_A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_output450_A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_output451_A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_output452_A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_output453_A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_output454_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_output455_A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_output456_A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_output457_A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_output458_A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_output459_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_output460_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_output461_A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_output468_A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_output481_A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_output483_A (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_output485_A (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_output486_A (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_output497_A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_output518_A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_output522_A (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_output523_A (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_output524_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_output525_A (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_output526_A (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_output527_A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_output528_A (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_output529_A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_output530_A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_output531_A (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_output532_A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_output533_A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_output536_A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A_N (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_output538_A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_output540_A (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_output541_A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_output542_A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_output543_A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_output544_A (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_output547_A (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_output548_A (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_output555_A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_output556_A (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_output557_A (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_output558_A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_output559_A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_output560_A (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_output561_A (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_output562_A (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__A1 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_output626_A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_output627_A (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_output628_A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_output629_A (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_output630_A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_output631_A (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_output633_A (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_output634_A (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_output635_A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_output636_A (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_output637_A (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA_output638_A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_output639_A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_output640_A (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_output664_A (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__A (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__A (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__A1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__B1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__S (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__S (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__S (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__A (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__A (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_output671_A (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_output672_A (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_output673_A (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_output674_A (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA_output675_A (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA_output677_A (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA_output678_A (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_output679_A (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_output680_A (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__7455__A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__7418__A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__7378__A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__CLK (.DIODE(clknet_leaf_1_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__CLK (.DIODE(clknet_leaf_1_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__CLK (.DIODE(clknet_leaf_1_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7311__CLK (.DIODE(clknet_leaf_2_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__CLK (.DIODE(clknet_leaf_2_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__CLK (.DIODE(clknet_leaf_2_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__CLK (.DIODE(clknet_leaf_2_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__CLK (.DIODE(clknet_leaf_2_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__CLK (.DIODE(clknet_leaf_2_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__CLK (.DIODE(clknet_leaf_2_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__CLK (.DIODE(clknet_leaf_4_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7018__CLK (.DIODE(clknet_leaf_4_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__CLK (.DIODE(clknet_leaf_4_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__CLK (.DIODE(clknet_leaf_4_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7168__CLK (.DIODE(clknet_leaf_4_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__CLK (.DIODE(clknet_leaf_4_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__CLK (.DIODE(clknet_leaf_4_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__CLK (.DIODE(clknet_leaf_4_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__CLK (.DIODE(clknet_leaf_4_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__CLK (.DIODE(clknet_leaf_5_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__CLK (.DIODE(clknet_leaf_5_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__CLK (.DIODE(clknet_leaf_5_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__CLK (.DIODE(clknet_leaf_5_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__CLK (.DIODE(clknet_leaf_5_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__CLK (.DIODE(clknet_leaf_7_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__CLK (.DIODE(clknet_leaf_7_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__CLK (.DIODE(clknet_leaf_7_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6984__CLK (.DIODE(clknet_leaf_7_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__CLK (.DIODE(clknet_leaf_7_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__CLK (.DIODE(clknet_leaf_7_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__CLK (.DIODE(clknet_leaf_7_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__CLK (.DIODE(clknet_leaf_7_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__CLK (.DIODE(clknet_leaf_7_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__CLK (.DIODE(clknet_leaf_9_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__CLK (.DIODE(clknet_leaf_9_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__CLK (.DIODE(clknet_leaf_9_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__CLK (.DIODE(clknet_leaf_9_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__CLK (.DIODE(clknet_leaf_9_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__CLK (.DIODE(clknet_leaf_9_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__CLK (.DIODE(clknet_leaf_9_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__CLK (.DIODE(clknet_leaf_9_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__CLK (.DIODE(clknet_leaf_9_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__CLK (.DIODE(clknet_leaf_9_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__CLK (.DIODE(clknet_leaf_10_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__CLK (.DIODE(clknet_leaf_10_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__CLK (.DIODE(clknet_leaf_10_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__CLK (.DIODE(clknet_leaf_10_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__CLK (.DIODE(clknet_leaf_10_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__CLK (.DIODE(clknet_leaf_10_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__CLK (.DIODE(clknet_leaf_10_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__CLK (.DIODE(clknet_leaf_10_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__CLK (.DIODE(clknet_leaf_10_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__CLK (.DIODE(clknet_leaf_10_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__CLK (.DIODE(clknet_leaf_11_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__CLK (.DIODE(clknet_leaf_11_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__CLK (.DIODE(clknet_leaf_11_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__CLK (.DIODE(clknet_leaf_11_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__CLK (.DIODE(clknet_leaf_11_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__CLK (.DIODE(clknet_leaf_11_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__CLK (.DIODE(clknet_leaf_11_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__CLK (.DIODE(clknet_leaf_11_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__CLK (.DIODE(clknet_leaf_11_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__CLK (.DIODE(clknet_leaf_11_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__CLK (.DIODE(clknet_leaf_12_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__CLK (.DIODE(clknet_leaf_12_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__CLK (.DIODE(clknet_leaf_12_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__CLK (.DIODE(clknet_leaf_12_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__CLK (.DIODE(clknet_leaf_12_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__CLK (.DIODE(clknet_leaf_12_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7173__CLK (.DIODE(clknet_leaf_12_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__CLK (.DIODE(clknet_leaf_13_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7121__CLK (.DIODE(clknet_leaf_13_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__CLK (.DIODE(clknet_leaf_13_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7136__CLK (.DIODE(clknet_leaf_13_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7185__CLK (.DIODE(clknet_leaf_13_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__CLK (.DIODE(clknet_leaf_13_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__CLK (.DIODE(clknet_leaf_13_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__CLK (.DIODE(clknet_leaf_13_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__CLK (.DIODE(clknet_leaf_13_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__CLK (.DIODE(clknet_leaf_13_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7309__CLK (.DIODE(clknet_leaf_19_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7251__CLK (.DIODE(clknet_leaf_19_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7264__CLK (.DIODE(clknet_leaf_19_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7307__CLK (.DIODE(clknet_leaf_19_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7308__CLK (.DIODE(clknet_leaf_19_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7379__A (.DIODE(clknet_leaf_19_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7200__CLK (.DIODE(clknet_leaf_22_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__CLK (.DIODE(clknet_leaf_22_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7203__CLK (.DIODE(clknet_leaf_22_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__CLK (.DIODE(clknet_leaf_22_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7229__CLK (.DIODE(clknet_leaf_22_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__CLK (.DIODE(clknet_leaf_22_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__CLK (.DIODE(clknet_leaf_22_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7276__CLK (.DIODE(clknet_leaf_22_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7271__CLK (.DIODE(clknet_leaf_25_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7260__CLK (.DIODE(clknet_leaf_25_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7258__CLK (.DIODE(clknet_leaf_25_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7259__CLK (.DIODE(clknet_leaf_25_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7270__CLK (.DIODE(clknet_leaf_25_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7283__CLK (.DIODE(clknet_leaf_25_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7262__CLK (.DIODE(clknet_leaf_25_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__CLK (.DIODE(clknet_leaf_25_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7233__CLK (.DIODE(clknet_leaf_26_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7234__CLK (.DIODE(clknet_leaf_26_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7273__CLK (.DIODE(clknet_leaf_26_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7247__CLK (.DIODE(clknet_leaf_26_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7246__CLK (.DIODE(clknet_leaf_26_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7245__CLK (.DIODE(clknet_leaf_26_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__CLK (.DIODE(clknet_leaf_26_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7284__CLK (.DIODE(clknet_leaf_26_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7286__CLK (.DIODE(clknet_leaf_26_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7285__CLK (.DIODE(clknet_leaf_26_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__CLK (.DIODE(clknet_leaf_27_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__CLK (.DIODE(clknet_leaf_27_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__CLK (.DIODE(clknet_leaf_27_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7192__CLK (.DIODE(clknet_leaf_27_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7194__CLK (.DIODE(clknet_leaf_27_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__CLK (.DIODE(clknet_leaf_27_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__CLK (.DIODE(clknet_leaf_27_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__CLK (.DIODE(clknet_leaf_27_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__CLK (.DIODE(clknet_leaf_27_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7232__CLK (.DIODE(clknet_leaf_27_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7208__CLK (.DIODE(clknet_leaf_27_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__CLK (.DIODE(clknet_leaf_28_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__CLK (.DIODE(clknet_leaf_28_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__CLK (.DIODE(clknet_leaf_28_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__CLK (.DIODE(clknet_leaf_28_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__CLK (.DIODE(clknet_leaf_28_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7187__CLK (.DIODE(clknet_leaf_28_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__CLK (.DIODE(clknet_leaf_28_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7217__CLK (.DIODE(clknet_leaf_28_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7191__CLK (.DIODE(clknet_leaf_28_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7218__CLK (.DIODE(clknet_leaf_28_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__CLK (.DIODE(clknet_leaf_28_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__CLK (.DIODE(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__CLK (.DIODE(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__CLK (.DIODE(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__CLK (.DIODE(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__CLK (.DIODE(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__CLK (.DIODE(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__CLK (.DIODE(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__CLK (.DIODE(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7128__CLK (.DIODE(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__CLK (.DIODE(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__CLK (.DIODE(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__CLK (.DIODE(clknet_leaf_29_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__CLK (.DIODE(clknet_leaf_30_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7102__CLK (.DIODE(clknet_leaf_30_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__CLK (.DIODE(clknet_leaf_30_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__CLK (.DIODE(clknet_leaf_30_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__CLK (.DIODE(clknet_leaf_30_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__CLK (.DIODE(clknet_leaf_30_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7155__CLK (.DIODE(clknet_leaf_30_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__CLK (.DIODE(clknet_leaf_30_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__CLK (.DIODE(clknet_leaf_30_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7153__CLK (.DIODE(clknet_leaf_30_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__CLK (.DIODE(clknet_leaf_32_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7109__CLK (.DIODE(clknet_leaf_32_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__CLK (.DIODE(clknet_leaf_32_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7093__CLK (.DIODE(clknet_leaf_32_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__CLK (.DIODE(clknet_leaf_32_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__CLK (.DIODE(clknet_leaf_32_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__CLK (.DIODE(clknet_leaf_32_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__CLK (.DIODE(clknet_leaf_32_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__CLK (.DIODE(clknet_leaf_32_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__CLK (.DIODE(clknet_leaf_32_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__CLK (.DIODE(clknet_leaf_32_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7139__CLK (.DIODE(clknet_leaf_33_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__CLK (.DIODE(clknet_leaf_33_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__CLK (.DIODE(clknet_leaf_33_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__CLK (.DIODE(clknet_leaf_33_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7152__CLK (.DIODE(clknet_leaf_33_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__CLK (.DIODE(clknet_leaf_33_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7179__CLK (.DIODE(clknet_leaf_33_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__CLK (.DIODE(clknet_leaf_33_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__CLK (.DIODE(clknet_leaf_33_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7171__CLK (.DIODE(clknet_leaf_33_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__CLK (.DIODE(clknet_leaf_34_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__CLK (.DIODE(clknet_leaf_34_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__CLK (.DIODE(clknet_leaf_34_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7148__CLK (.DIODE(clknet_leaf_34_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__CLK (.DIODE(clknet_leaf_34_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__CLK (.DIODE(clknet_leaf_34_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__CLK (.DIODE(clknet_leaf_34_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__CLK (.DIODE(clknet_leaf_34_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7098__CLK (.DIODE(clknet_leaf_35_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__CLK (.DIODE(clknet_leaf_35_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7174__CLK (.DIODE(clknet_leaf_35_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__CLK (.DIODE(clknet_leaf_35_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__CLK (.DIODE(clknet_leaf_35_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__CLK (.DIODE(clknet_leaf_35_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7170__CLK (.DIODE(clknet_leaf_35_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__CLK (.DIODE(clknet_leaf_35_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7147__CLK (.DIODE(clknet_leaf_35_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__CLK (.DIODE(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__CLK (.DIODE(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__CLK (.DIODE(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__CLK (.DIODE(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__CLK (.DIODE(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__CLK (.DIODE(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__CLK (.DIODE(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__CLK (.DIODE(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__CLK (.DIODE(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__CLK (.DIODE(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__CLK (.DIODE(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__CLK (.DIODE(clknet_leaf_36_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__CLK (.DIODE(clknet_leaf_37_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__CLK (.DIODE(clknet_leaf_37_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__CLK (.DIODE(clknet_leaf_37_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__CLK (.DIODE(clknet_leaf_37_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7048__CLK (.DIODE(clknet_leaf_37_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__CLK (.DIODE(clknet_leaf_37_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__CLK (.DIODE(clknet_leaf_37_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__CLK (.DIODE(clknet_leaf_37_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__CLK (.DIODE(clknet_leaf_37_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__CLK (.DIODE(clknet_leaf_38_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__CLK (.DIODE(clknet_leaf_38_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__CLK (.DIODE(clknet_leaf_38_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__CLK (.DIODE(clknet_leaf_38_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__CLK (.DIODE(clknet_leaf_38_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__CLK (.DIODE(clknet_leaf_38_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__CLK (.DIODE(clknet_leaf_39_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__CLK (.DIODE(clknet_leaf_39_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__CLK (.DIODE(clknet_leaf_39_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__CLK (.DIODE(clknet_leaf_39_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__CLK (.DIODE(clknet_leaf_39_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__CLK (.DIODE(clknet_leaf_39_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__CLK (.DIODE(clknet_leaf_39_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__CLK (.DIODE(clknet_leaf_39_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__CLK (.DIODE(clknet_leaf_41_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__CLK (.DIODE(clknet_leaf_41_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__CLK (.DIODE(clknet_leaf_41_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__CLK (.DIODE(clknet_leaf_41_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__CLK (.DIODE(clknet_leaf_41_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__CLK (.DIODE(clknet_leaf_41_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__CLK (.DIODE(clknet_leaf_41_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__CLK (.DIODE(clknet_leaf_41_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__CLK (.DIODE(clknet_leaf_41_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__CLK (.DIODE(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__CLK (.DIODE(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__CLK (.DIODE(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__CLK (.DIODE(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__CLK (.DIODE(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__CLK (.DIODE(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__CLK (.DIODE(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__CLK (.DIODE(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__CLK (.DIODE(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__CLK (.DIODE(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__CLK (.DIODE(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__CLK (.DIODE(clknet_leaf_42_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7297__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7298__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7293__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7294__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7292__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__CLK (.DIODE(clknet_leaf_43_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__CLK (.DIODE(clknet_leaf_44_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7296__CLK (.DIODE(clknet_leaf_44_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7299__CLK (.DIODE(clknet_leaf_44_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7300__CLK (.DIODE(clknet_leaf_44_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7295__CLK (.DIODE(clknet_leaf_44_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7291__CLK (.DIODE(clknet_leaf_44_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__CLK (.DIODE(clknet_leaf_44_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7301__CLK (.DIODE(clknet_leaf_44_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__CLK (.DIODE(clknet_leaf_44_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__CLK (.DIODE(clknet_leaf_44_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__CLK (.DIODE(clknet_leaf_44_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__CLK (.DIODE(clknet_leaf_45_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__CLK (.DIODE(clknet_leaf_46_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__CLK (.DIODE(clknet_leaf_46_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__CLK (.DIODE(clknet_leaf_46_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__CLK (.DIODE(clknet_leaf_46_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__CLK (.DIODE(clknet_leaf_46_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__CLK (.DIODE(clknet_leaf_46_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__CLK (.DIODE(clknet_leaf_46_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__CLK (.DIODE(clknet_leaf_46_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__CLK (.DIODE(clknet_leaf_48_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__CLK (.DIODE(clknet_leaf_48_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__CLK (.DIODE(clknet_leaf_48_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__CLK (.DIODE(clknet_leaf_48_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__CLK (.DIODE(clknet_leaf_48_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__CLK (.DIODE(clknet_leaf_48_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__CLK (.DIODE(clknet_leaf_48_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__CLK (.DIODE(clknet_leaf_48_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__CLK (.DIODE(clknet_leaf_49_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__CLK (.DIODE(clknet_leaf_50_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__CLK (.DIODE(clknet_leaf_50_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__CLK (.DIODE(clknet_leaf_50_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__CLK (.DIODE(clknet_leaf_50_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__CLK (.DIODE(clknet_leaf_50_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__CLK (.DIODE(clknet_leaf_50_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__CLK (.DIODE(clknet_leaf_50_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__CLK (.DIODE(clknet_leaf_50_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__CLK (.DIODE(clknet_leaf_50_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__CLK (.DIODE(clknet_leaf_53_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__CLK (.DIODE(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__CLK (.DIODE(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__CLK (.DIODE(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__CLK (.DIODE(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__CLK (.DIODE(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__CLK (.DIODE(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__CLK (.DIODE(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__CLK (.DIODE(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__CLK (.DIODE(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__CLK (.DIODE(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__CLK (.DIODE(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__CLK (.DIODE(clknet_leaf_54_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__CLK (.DIODE(clknet_leaf_56_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__CLK (.DIODE(clknet_leaf_57_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__CLK (.DIODE(clknet_leaf_57_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__CLK (.DIODE(clknet_leaf_57_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__CLK (.DIODE(clknet_leaf_57_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__CLK (.DIODE(clknet_leaf_57_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__CLK (.DIODE(clknet_leaf_57_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__CLK (.DIODE(clknet_leaf_57_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__CLK (.DIODE(clknet_leaf_58_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__CLK (.DIODE(clknet_leaf_58_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__CLK (.DIODE(clknet_leaf_58_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__CLK (.DIODE(clknet_leaf_58_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__CLK (.DIODE(clknet_leaf_58_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__CLK (.DIODE(clknet_leaf_58_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__CLK (.DIODE(clknet_leaf_58_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__CLK (.DIODE(clknet_leaf_58_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__CLK (.DIODE(clknet_leaf_58_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__CLK (.DIODE(clknet_leaf_59_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__CLK (.DIODE(clknet_leaf_59_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__CLK (.DIODE(clknet_leaf_59_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__CLK (.DIODE(clknet_leaf_59_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__CLK (.DIODE(clknet_leaf_59_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__CLK (.DIODE(clknet_leaf_59_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__CLK (.DIODE(clknet_leaf_59_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__CLK (.DIODE(clknet_leaf_59_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__CLK (.DIODE(clknet_leaf_59_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__CLK (.DIODE(clknet_leaf_59_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__CLK (.DIODE(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__CLK (.DIODE(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__CLK (.DIODE(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__CLK (.DIODE(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7302__CLK (.DIODE(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__CLK (.DIODE(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__CLK (.DIODE(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__CLK (.DIODE(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__CLK (.DIODE(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__CLK (.DIODE(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__CLK (.DIODE(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__CLK (.DIODE(clknet_leaf_62_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__CLK (.DIODE(clknet_leaf_63_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__CLK (.DIODE(clknet_leaf_63_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__CLK (.DIODE(clknet_leaf_63_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__CLK (.DIODE(clknet_leaf_63_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__CLK (.DIODE(clknet_leaf_63_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__CLK (.DIODE(clknet_leaf_63_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__CLK (.DIODE(clknet_leaf_63_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__CLK (.DIODE(clknet_leaf_63_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__CLK (.DIODE(clknet_leaf_63_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__CLK (.DIODE(clknet_leaf_63_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__CLK (.DIODE(clknet_leaf_66_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__CLK (.DIODE(clknet_leaf_68_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6842__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6846__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__CLK (.DIODE(clknet_leaf_69_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__CLK (.DIODE(clknet_leaf_70_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__CLK (.DIODE(clknet_leaf_70_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__CLK (.DIODE(clknet_leaf_70_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__CLK (.DIODE(clknet_leaf_70_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__CLK (.DIODE(clknet_leaf_70_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__CLK (.DIODE(clknet_leaf_70_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__CLK (.DIODE(clknet_leaf_70_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__CLK (.DIODE(clknet_leaf_70_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__CLK (.DIODE(clknet_leaf_70_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__CLK (.DIODE(clknet_leaf_70_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__CLK (.DIODE(clknet_leaf_70_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6881__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__CLK (.DIODE(clknet_leaf_71_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__CLK (.DIODE(clknet_leaf_75_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__CLK (.DIODE(clknet_leaf_75_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__CLK (.DIODE(clknet_leaf_75_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__CLK (.DIODE(clknet_leaf_75_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__CLK (.DIODE(clknet_leaf_75_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__CLK (.DIODE(clknet_leaf_75_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__CLK (.DIODE(clknet_leaf_75_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6926__CLK (.DIODE(clknet_leaf_76_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__CLK (.DIODE(clknet_leaf_76_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__CLK (.DIODE(clknet_leaf_76_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__CLK (.DIODE(clknet_leaf_76_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__CLK (.DIODE(clknet_leaf_76_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__CLK (.DIODE(clknet_leaf_76_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__CLK (.DIODE(clknet_leaf_76_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__CLK (.DIODE(clknet_leaf_76_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__CLK (.DIODE(clknet_leaf_76_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__CLK (.DIODE(clknet_leaf_76_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__CLK (.DIODE(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__CLK (.DIODE(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__CLK (.DIODE(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__CLK (.DIODE(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__CLK (.DIODE(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__CLK (.DIODE(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__CLK (.DIODE(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__CLK (.DIODE(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__CLK (.DIODE(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__CLK (.DIODE(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7074__CLK (.DIODE(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__CLK (.DIODE(clknet_leaf_79_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__CLK (.DIODE(clknet_leaf_80_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__CLK (.DIODE(clknet_leaf_80_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__CLK (.DIODE(clknet_leaf_80_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__CLK (.DIODE(clknet_leaf_80_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7061__CLK (.DIODE(clknet_leaf_80_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__CLK (.DIODE(clknet_leaf_80_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__CLK (.DIODE(clknet_leaf_80_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__CLK (.DIODE(clknet_leaf_80_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__CLK (.DIODE(clknet_leaf_80_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7058__CLK (.DIODE(clknet_leaf_80_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__CLK (.DIODE(clknet_leaf_80_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__CLK (.DIODE(clknet_leaf_81_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__CLK (.DIODE(clknet_leaf_81_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__CLK (.DIODE(clknet_leaf_81_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__CLK (.DIODE(clknet_leaf_81_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__CLK (.DIODE(clknet_leaf_81_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__CLK (.DIODE(clknet_leaf_81_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__CLK (.DIODE(clknet_leaf_81_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7019__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__CLK (.DIODE(clknet_leaf_82_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__CLK (.DIODE(clknet_leaf_85_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6958__CLK (.DIODE(clknet_leaf_85_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__CLK (.DIODE(clknet_leaf_85_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__CLK (.DIODE(clknet_leaf_85_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__CLK (.DIODE(clknet_leaf_85_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__CLK (.DIODE(clknet_leaf_85_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__CLK (.DIODE(clknet_leaf_85_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__CLK (.DIODE(clknet_leaf_85_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__CLK (.DIODE(clknet_leaf_85_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__CLK (.DIODE(clknet_leaf_85_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__CLK (.DIODE(clknet_leaf_85_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__CLK (.DIODE(clknet_leaf_86_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__CLK (.DIODE(clknet_leaf_86_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__CLK (.DIODE(clknet_leaf_86_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__CLK (.DIODE(clknet_leaf_86_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__CLK (.DIODE(clknet_leaf_86_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__CLK (.DIODE(clknet_leaf_86_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__CLK (.DIODE(clknet_leaf_86_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7341__A (.DIODE(clknet_leaf_92_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7290__CLK (.DIODE(clknet_leaf_92_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7417__A (.DIODE(clknet_leaf_92_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__CLK (.DIODE(clknet_leaf_93_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__CLK (.DIODE(clknet_leaf_93_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7287__CLK (.DIODE(clknet_leaf_93_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7289__CLK (.DIODE(clknet_leaf_93_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7085__CLK (.DIODE(clknet_leaf_93_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__CLK (.DIODE(clknet_leaf_93_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__CLK (.DIODE(clknet_leaf_93_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_core_clock_A (.DIODE(clknet_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_core_clock_A (.DIODE(clknet_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_core_clock_A (.DIODE(clknet_1_0_1_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_core_clock_A (.DIODE(clknet_1_0_1_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_core_clock_A (.DIODE(clknet_1_1_1_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_core_clock_A (.DIODE(clknet_1_1_1_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_core_clock_A (.DIODE(clknet_2_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_core_clock_A (.DIODE(clknet_2_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_core_clock_A (.DIODE(clknet_2_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_core_clock_A (.DIODE(clknet_2_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_core_clock_A (.DIODE(clknet_2_2_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_core_clock_A (.DIODE(clknet_2_2_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_core_clock_A (.DIODE(clknet_2_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_core_clock_A (.DIODE(clknet_2_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_core_clock_A (.DIODE(clknet_3_0_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_core_clock_A (.DIODE(clknet_3_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_core_clock_A (.DIODE(clknet_3_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_core_clock_A (.DIODE(clknet_3_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_core_clock_A (.DIODE(clknet_3_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_core_clock_A (.DIODE(clknet_3_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_core_clock_A (.DIODE(clknet_3_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_core_clock_A (.DIODE(clknet_3_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_core_clock_A (.DIODE(clknet_3_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_core_clock_A (.DIODE(clknet_3_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_core_clock_A (.DIODE(clknet_3_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_core_clock_A (.DIODE(clknet_3_1_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_core_clock_A (.DIODE(clknet_3_2_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_core_clock_A (.DIODE(clknet_3_2_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_core_clock_A (.DIODE(clknet_3_2_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_core_clock_A (.DIODE(clknet_3_2_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_core_clock_A (.DIODE(clknet_3_2_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_core_clock_A (.DIODE(clknet_3_2_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_core_clock_A (.DIODE(clknet_3_2_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_core_clock_A (.DIODE(clknet_3_2_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_1_0_core_clock_A (.DIODE(clknet_3_2_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__CLK (.DIODE(clknet_3_2_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_core_clock_A (.DIODE(clknet_3_3_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_core_clock_A (.DIODE(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_core_clock_A (.DIODE(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_core_clock_A (.DIODE(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_core_clock_A (.DIODE(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_core_clock_A (.DIODE(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_core_clock_A (.DIODE(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_core_clock_A (.DIODE(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_core_clock_A (.DIODE(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_core_clock_A (.DIODE(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_core_clock_A (.DIODE(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_core_clock_A (.DIODE(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_core_clock_A (.DIODE(clknet_3_4_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_core_clock_A (.DIODE(clknet_3_5_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_core_clock_A (.DIODE(clknet_3_5_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_core_clock_A (.DIODE(clknet_3_5_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_core_clock_A (.DIODE(clknet_3_5_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_core_clock_A (.DIODE(clknet_3_5_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_core_clock_A (.DIODE(clknet_3_5_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_core_clock_A (.DIODE(clknet_3_5_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_core_clock_A (.DIODE(clknet_3_5_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_core_clock_A (.DIODE(clknet_3_5_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_core_clock_A (.DIODE(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_core_clock_A (.DIODE(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_core_clock_A (.DIODE(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_core_clock_A (.DIODE(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_2_0_core_clock_A (.DIODE(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_core_clock_A (.DIODE(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_core_clock_A (.DIODE(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_core_clock_A (.DIODE(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_core_clock_A (.DIODE(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_core_clock_A (.DIODE(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_core_clock_A (.DIODE(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_core_clock_A (.DIODE(clknet_3_6_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_core_clock_A (.DIODE(clknet_3_7_0_core_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__7435__A (.DIODE(clknet_opt_1_0_core_clock));
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_623 ();
 assign c0_i_core_int_sreg[10] = net719;
 assign c0_i_core_int_sreg[11] = net720;
 assign c0_i_core_int_sreg[12] = net721;
 assign c0_i_core_int_sreg[13] = net722;
 assign c0_i_core_int_sreg[14] = net723;
 assign c0_i_core_int_sreg[15] = net724;
 assign c0_i_core_int_sreg[2] = net711;
 assign c0_i_core_int_sreg[3] = net712;
 assign c0_i_core_int_sreg[4] = net713;
 assign c0_i_core_int_sreg[5] = net714;
 assign c0_i_core_int_sreg[6] = net715;
 assign c0_i_core_int_sreg[7] = net716;
 assign c0_i_core_int_sreg[8] = net717;
 assign c0_i_core_int_sreg[9] = net718;
 assign c1_i_core_int_sreg[10] = net733;
 assign c1_i_core_int_sreg[11] = net734;
 assign c1_i_core_int_sreg[12] = net735;
 assign c1_i_core_int_sreg[13] = net736;
 assign c1_i_core_int_sreg[14] = net737;
 assign c1_i_core_int_sreg[15] = net738;
 assign c1_i_core_int_sreg[2] = net725;
 assign c1_i_core_int_sreg[3] = net726;
 assign c1_i_core_int_sreg[4] = net727;
 assign c1_i_core_int_sreg[5] = net728;
 assign c1_i_core_int_sreg[6] = net729;
 assign c1_i_core_int_sreg[7] = net730;
 assign c1_i_core_int_sreg[8] = net731;
 assign c1_i_core_int_sreg[9] = net732;
 assign c1_i_irq = net739;
endmodule

