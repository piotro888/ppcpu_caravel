magic
tech sky130B
magscale 1 2
timestamp 1662739868
<< nwell >>
rect 1066 37253 38862 37574
rect 1066 36165 38862 36731
rect 1066 35077 38862 35643
rect 1066 33989 38862 34555
rect 1066 32901 38862 33467
rect 1066 31813 38862 32379
rect 1066 30725 38862 31291
rect 1066 29637 38862 30203
rect 1066 28549 38862 29115
rect 1066 27461 38862 28027
rect 1066 26373 38862 26939
rect 1066 25285 38862 25851
rect 1066 24197 38862 24763
rect 1066 23109 38862 23675
rect 1066 22021 38862 22587
rect 1066 20933 38862 21499
rect 1066 19845 38862 20411
rect 1066 18757 38862 19323
rect 1066 17669 38862 18235
rect 1066 16581 38862 17147
rect 1066 15493 38862 16059
rect 1066 14405 38862 14971
rect 1066 13317 38862 13883
rect 1066 12229 38862 12795
rect 1066 11141 38862 11707
rect 1066 10053 38862 10619
rect 1066 8965 38862 9531
rect 1066 7877 38862 8443
rect 1066 6789 38862 7355
rect 1066 5701 38862 6267
rect 1066 4613 38862 5179
rect 1066 3525 38862 4091
rect 1066 2437 38862 3003
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 1104 2128 38824 37584
<< metal2 >>
rect 6642 39200 6698 40000
rect 19982 39200 20038 40000
rect 33322 39200 33378 40000
<< obsm2 >>
rect 4214 39144 6586 39200
rect 6754 39144 19926 39200
rect 20094 39144 33266 39200
rect 33434 39144 35242 39200
rect 4214 2139 35242 39144
<< obsm3 >>
rect 4210 2143 35246 37569
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal2 s 6642 39200 6698 40000 6 a
port 1 nsew signal input
rlabel metal2 s 19982 39200 20038 40000 6 b
port 2 nsew signal input
rlabel metal2 s 33322 39200 33378 40000 6 c
port 3 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 4 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 4 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 414446
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/t2/runs/22_09_09_18_10/results/signoff/t2.magic.gds
string GDS_START 37058
<< end >>

