* NGSPICE file created from RAM32.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlclkp_1 abstract view
.subckt sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

.subckt RAM32 A0[0] A0[1] A0[2] A0[3] A0[4] CLK Di0[0] Di0[10] Di0[11] Di0[12] Di0[13]
+ Di0[14] Di0[15] Di0[16] Di0[17] Di0[18] Di0[19] Di0[1] Di0[20] Di0[21] Di0[22] Di0[23]
+ Di0[24] Di0[25] Di0[26] Di0[27] Di0[28] Di0[29] Di0[2] Di0[30] Di0[31] Di0[32] Di0[33]
+ Di0[34] Di0[35] Di0[36] Di0[37] Di0[38] Di0[39] Di0[3] Di0[40] Di0[41] Di0[42] Di0[43]
+ Di0[44] Di0[45] Di0[46] Di0[47] Di0[48] Di0[49] Di0[4] Di0[50] Di0[51] Di0[52] Di0[53]
+ Di0[54] Di0[55] Di0[56] Di0[57] Di0[58] Di0[59] Di0[5] Di0[60] Di0[61] Di0[62] Di0[63]
+ Di0[6] Di0[7] Di0[8] Di0[9] Do0[0] Do0[10] Do0[11] Do0[12] Do0[13] Do0[14] Do0[15]
+ Do0[16] Do0[17] Do0[18] Do0[19] Do0[1] Do0[20] Do0[21] Do0[22] Do0[23] Do0[24] Do0[25]
+ Do0[26] Do0[27] Do0[28] Do0[29] Do0[2] Do0[30] Do0[31] Do0[32] Do0[33] Do0[34] Do0[35]
+ Do0[36] Do0[37] Do0[38] Do0[39] Do0[3] Do0[40] Do0[41] Do0[42] Do0[43] Do0[44] Do0[45]
+ Do0[46] Do0[47] Do0[48] Do0[49] Do0[4] Do0[50] Do0[51] Do0[52] Do0[53] Do0[54] Do0[55]
+ Do0[56] Do0[57] Do0[58] Do0[59] Do0[5] Do0[60] Do0[61] Do0[62] Do0[63] Do0[6] Do0[7]
+ Do0[8] Do0[9] EN0 VGND VPWR WE0[0] WE0[1] WE0[2] WE0[3] WE0[4] WE0[5] WE0[6] WE0[7]
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG net80 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_39_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV_81 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_62_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[44\].__cell__ Di0[44] VGND VGND VPWR VPWR DIBUF\[44\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_132_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CLKINV_55 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__inv_1
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WEBUF\[5\].__cell__ SLICE\[0\].RAM8.WEBUF\[5\].A VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WEBUF\[5\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_54_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_123_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_76_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG net27 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_9_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_86_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_28_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[2\] Do0_REG.CLKBUF\[7\] BYTE\[7\].FLOATBUF0\[58\].Z
+ VGND VGND VPWR VPWR Do0[58] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CLKINV_103 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_128_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG net184 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_117_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_104_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_120_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_19_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG net140 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WEBUF\[7\].__cell__ SLICE\[0\].RAM8.WEBUF\[7\].A VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WEBUF\[7\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_101_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[2\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_3_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CLKINV_87 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__inv_1
XFILLER_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CLKINV_135 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__inv_1
XFILLER_48_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV_99 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__inv_1
XFILLER_74_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV_162 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__inv_1
XFILLER_15_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CLKINV_192 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_128_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_127_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_97_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG net244 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[6\] Do0_REG.CLKBUF\[3\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VGND VGND VPWR VPWR Do0[30] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_87_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_79_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_39_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV_194 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__inv_1
XFILLER_85_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[7\].FLOATBUF0\[59\].__cell__ BYTE\[7\].FLOATBUF0\[56\].A BYTE\[7\].FLOATBUF0\[56\].TE_B
+ VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_71_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CLKINV_63 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_107_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.DEC0.AND4 SLICE\[1\].RAM8.DEC0.A_buf\[0\] SLICE\[1\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[4\].W.SEL0 sky130_fd_sc_hd__and4bb_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG net38 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_106_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XBYTE\[3\].FLOATBUF0\[27\].__cell__ BYTE\[3\].FLOATBUF0\[24\].A BYTE\[3\].FLOATBUF0\[24\].TE_B
+ VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_48_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_63_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_112_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[34\].__cell__ Di0[34] VGND VGND VPWR VPWR DIBUF\[34\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_50_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_106_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG net151 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_53_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_103_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[6\].FLOATBUF0\[50\].__cell__ BYTE\[6\].FLOATBUF0\[48\].A BYTE\[6\].FLOATBUF0\[48\].TE_B
+ VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_32_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_132_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_27_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG net98 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_117_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_58_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_73_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CLKINV_95 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__inv_1
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG net255 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_5_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG net211 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_99_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_67_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_94_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[1\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV_164 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__inv_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_88_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_73_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_127_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_6_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_111_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_84_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_49_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV_249 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[3\] Do0_REG.CLKBUF\[0\] BYTE\[0\].FLOATBUF0\[3\].Z
+ VGND VGND VPWR VPWR Do0[3] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG net5 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_114_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_128_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_128_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.DEC0.ENBUF SLICE\[0\].RAM8.DEC0.EN VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.EN_buf
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_109_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_66_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV_196 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_128_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_119_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CLKINV_230 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_88_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_70_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG net109 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_47_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDIBUF\[24\].__cell__ Di0[24] VGND VGND VPWR VPWR DIBUF\[24\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG net65 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_116_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_69_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[63\].__cell__ Di0[63] VGND VGND VPWR VPWR DIBUF\[63\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_119_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.DEC0.AND5 SLICE\[1\].RAM8.DEC0.A_buf\[1\] SLICE\[1\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[5\].W.SEL0 sky130_fd_sc_hd__and4b_2
XFILLER_107_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_96_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG net222 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[2\].FLOATBUF0\[19\].__cell__ BYTE\[2\].FLOATBUF0\[16\].A BYTE\[2\].FLOATBUF0\[16\].TE_B
+ VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_4_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_131_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_81_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG net169 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_13_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_126_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[8\].__cell__ Di0[8] VGND VGND VPWR VPWR DIBUF\[8\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG net16 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_122_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_32_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[3\] Do0_REG.CLKBUF\[5\] BYTE\[5\].FLOATBUF0\[43\].Z
+ VGND VGND VPWR VPWR Do0[43] sky130_fd_sc_hd__dfxtp_1
XBYTE\[5\].FLOATBUF0\[42\].__cell__ BYTE\[5\].FLOATBUF0\[40\].A BYTE\[5\].FLOATBUF0\[40\].TE_B
+ VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CLKINV_166 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__inv_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[1\].FLOATBUF0\[10\].__cell__ BYTE\[1\].FLOATBUF0\[10\].A BYTE\[1\].FLOATBUF0\[10\].TE_B
+ VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_23_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[0\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_109_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_14_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XWEBUF\[4\].__cell__ WE0[4] VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[4\].A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_107_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_110_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_1_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_45_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_60_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG net120 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CLKINV_198 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG net76 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_132_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_85_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[7\] Do0_REG.CLKBUF\[1\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VGND VGND VPWR VPWR Do0[15] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV_202 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__inv_1
XFILLER_110_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CLKINV_232 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__inv_1
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_114_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_117_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_74_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[14\].__cell__ Di0[14] VGND VGND VPWR VPWR DIBUF\[14\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG net180 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_10_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_127_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_97_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XDIBUF\[53\].__cell__ Di0[53] VGND VGND VPWR VPWR DIBUF\[53\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_65_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV_106 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__inv_1
XFILLER_52_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_71_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_8_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_3_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_120_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_97_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_53_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.CLKBUF.__cell__ CLKBUF.X VGND VGND VPWR VPWR SLICE\[2\].RAM8.CLKBUF.X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_21_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.DEC0.AND6 SLICE\[1\].RAM8.DEC0.A_buf\[0\] SLICE\[1\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[6\].W.SEL0 sky130_fd_sc_hd__and4b_2
XFILLER_106_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_121_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV_138 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__inv_1
XFILLER_130_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CLKINV_168 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__inv_1
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[0\] Do0_REG.CLKBUF\[2\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VGND VGND VPWR VPWR Do0[16] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_61_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG net87 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_106_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_67_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_62_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_30_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_116_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_116_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_85_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_107_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[7\] Do0_REG.CLKBUF\[6\] BYTE\[6\].FLOATBUF0\[55\].Z
+ VGND VGND VPWR VPWR Do0[55] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG net200 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG net34 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_4_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[4\].FLOATBUF0\[34\].__cell__ BYTE\[4\].FLOATBUF0\[32\].A BYTE\[4\].FLOATBUF0\[32\].TE_B
+ VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_35_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG net191 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_50_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_117_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_131_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV_204 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG net147 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_108_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WEBUF\[2\].__cell__ SLICE\[0\].RAM8.WEBUF\[2\].A VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WEBUF\[2\].X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_9_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_4_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[0\].FLOATBUF0\[7\].__cell__ BYTE\[0\].FLOATBUF0\[0\].A BYTE\[0\].FLOATBUF0\[0\].TE_B
+ VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_100_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_53_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV_108 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_52_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_118_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_96_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[43\].__cell__ Di0[43] VGND VGND VPWR VPWR DIBUF\[43\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_77_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG net251 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WEBUF\[4\].__cell__ SLICE\[0\].RAM8.WEBUF\[4\].A VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WEBUF\[4\].X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_68_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[0\] Do0_REG.CLKBUF\[7\] BYTE\[7\].FLOATBUF0\[56\].Z
+ VGND VGND VPWR VPWR Do0[56] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_124_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_59_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_100_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_111_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_65_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG net45 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_60_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_20_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV_12 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__inv_1
XFILLER_28_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG net1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WEBUF\[6\].__cell__ SLICE\[0\].RAM8.WEBUF\[6\].A VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WEBUF\[6\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_109_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_3_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_47_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG net158 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_116_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_111_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_65_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[4\] Do0_REG.CLKBUF\[3\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VGND VGND VPWR VPWR Do0[28] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.DEC0.AND7 SLICE\[1\].RAM8.DEC0.A_buf\[0\] SLICE\[1\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[7\].W.SEL0 sky130_fd_sc_hd__and4_2
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_130_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_91_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_29_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_71_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_8_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_121_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG net105 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CLKINV_206 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV_233 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_102_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.CLKBUF.__cell__ CLKBUF.X VGND VGND VPWR VPWR SLICE\[0\].RAM8.CLKBUF.X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_72_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG net218 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XBYTE\[7\].FLOATBUF0\[58\].__cell__ BYTE\[7\].FLOATBUF0\[56\].A BYTE\[7\].FLOATBUF0\[56\].TE_B
+ VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_4_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_94_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XBYTE\[3\].FLOATBUF0\[26\].__cell__ BYTE\[3\].FLOATBUF0\[24\].A BYTE\[3\].FLOATBUF0\[24\].TE_B
+ VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG net56 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_5_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[33\].__cell__ Di0[33] VGND VGND VPWR VPWR DIBUF\[33\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_122_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_67_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_1_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG net12 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_9_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_94_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_103_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_55_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_23_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV_20 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_132_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_104_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_77_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_10_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_127_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_6_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV_169 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_49_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_91_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_17_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG net116 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_82_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_63_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_59_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_128_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_89_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[1\] Do0_REG.CLKBUF\[0\] BYTE\[0\].FLOATBUF0\[1\].Z
+ VGND VGND VPWR VPWR Do0[1] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG net229 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_119_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CLKINV_150 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__inv_1
XFILLER_118_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[1\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_87_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_68_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_83_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_70_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_34_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_50_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CLKINV_208 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_105_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV_235 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__inv_1
XFILLER_75_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_62_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_7_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CLKINV_38 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_57_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG net23 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_112_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_130_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_12_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_39_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG net136 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_119_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XDIBUF\[23\].__cell__ Di0[23] VGND VGND VPWR VPWR DIBUF\[23\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_1_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_76_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_29_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG net127 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_56_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[62\].__cell__ Di0[62] VGND VGND VPWR VPWR DIBUF\[62\].X sky130_fd_sc_hd__clkbuf_16
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_39_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_63_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG net83 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_50_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XBYTE\[2\].FLOATBUF0\[18\].__cell__ BYTE\[2\].FLOATBUF0\[16\].A BYTE\[2\].FLOATBUF0\[16\].TE_B
+ VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_85_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CLKINV_120 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__inv_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG net240 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_60_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[1\] Do0_REG.CLKBUF\[5\] BYTE\[5\].FLOATBUF0\[41\].Z
+ VGND VGND VPWR VPWR Do0[41] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_9_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG net196 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_95_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[7\].__cell__ Di0[7] VGND VGND VPWR VPWR DIBUF\[7\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_82_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_90_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_109_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_105_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG net187 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[5\].FLOATBUF0\[41\].__cell__ BYTE\[5\].FLOATBUF0\[40\].A BYTE\[5\].FLOATBUF0\[40\].TE_B
+ VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_86_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_100_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_54_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_6_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CLKINV_152 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__inv_1
XFILLER_96_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_77_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CLKINV_46 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__inv_1
XFILLER_33_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV_58 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__inv_1
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_102_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XWEBUF\[3\].__cell__ WE0[3] VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[3\].A sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CLKINV_237 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__inv_1
XFILLER_24_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_3_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_30_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_97_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[5\] Do0_REG.CLKBUF\[1\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VGND VGND VPWR VPWR Do0[13] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_2_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_125_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_96_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG net94 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_117_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_93_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_86_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_74_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_62_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CLKINV_78 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_61_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_119_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_106_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG net207 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDIBUF\[13\].__cell__ Di0[13] VGND VGND VPWR VPWR DIBUF\[13\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG net41 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_45_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[52\].__cell__ Di0[52] VGND VGND VPWR VPWR DIBUF\[52\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_8_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_121_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_128_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG net154 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_80_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_107_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_103_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_72_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CLKINV_54 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__inv_1
XFILLER_39_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_54_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_53_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_42_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CLKINV_181 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__inv_1
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_107_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_123_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[5\] Do0_REG.CLKBUF\[6\] BYTE\[6\].FLOATBUF0\[53\].Z
+ VGND VGND VPWR VPWR Do0[53] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_123_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV_209 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__inv_1
XFILLER_60_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CLKINV_239 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__inv_1
XFILLER_9_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_95_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_51_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_50_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_117_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_85_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[4\].FLOATBUF0\[33\].__cell__ BYTE\[4\].FLOATBUF0\[32\].A BYTE\[4\].FLOATBUF0\[32\].TE_B
+ VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG net52 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_104_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.Do_CLKBUF\[7\] Do0_REG.CLK_buf VGND VGND VPWR VPWR Do0_REG.CLKBUF\[7\] sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_32_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_99_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CLKINV_86 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__inv_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV_98 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__inv_1
XFILLER_36_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_3_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_78_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WEBUF\[1\].__cell__ SLICE\[0\].RAM8.WEBUF\[1\].A VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WEBUF\[1\].X sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_120_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG net165 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_128_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_49_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[0\].FLOATBUF0\[6\].__cell__ BYTE\[0\].FLOATBUF0\[0\].A BYTE\[0\].FLOATBUF0\[0\].TE_B
+ VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_33_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_51_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDIBUF\[42\].__cell__ Di0[42] VGND VGND VPWR VPWR DIBUF\[42\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_79_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV_121 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__inv_1
XFILLER_87_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_115_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.DEC0.ENBUF SLICE\[3\].RAM8.DEC0.EN VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.EN_buf
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WEBUF\[3\].__cell__ SLICE\[0\].RAM8.WEBUF\[3\].A VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WEBUF\[3\].X sky130_fd_sc_hd__clkbuf_2
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_42_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CLKINV_62 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_130_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_106_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_130_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG net225 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_44_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.DEC0.ABUF\[1\] A0BUF\[1\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.A_buf\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_125_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG net72 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_15_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV_153 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__inv_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CLKINV_183 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__inv_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WEBUF\[5\].__cell__ SLICE\[0\].RAM8.WEBUF\[5\].A VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WEBUF\[5\].X sky130_fd_sc_hd__clkbuf_2
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CG net63 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_81_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_81_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_80_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[2\] Do0_REG.CLKBUF\[3\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VGND VGND VPWR VPWR Do0[26] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG net19 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_91_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_44_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_126_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_106_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_79_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_63_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG net176 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_90_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CLKINV_94 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__inv_1
XFILLER_117_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_89_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG net132 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WEBUF\[7\].__cell__ SLICE\[0\].RAM8.WEBUF\[7\].A VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WEBUF\[7\].X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_108_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_123_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_107_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_123_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_40_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG net123 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_51_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[7\].FLOATBUF0\[57\].__cell__ BYTE\[7\].FLOATBUF0\[56\].A BYTE\[7\].FLOATBUF0\[56\].TE_B
+ VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_85_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_42_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_10_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_127_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_123_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBYTE\[3\].FLOATBUF0\[25\].__cell__ BYTE\[3\].FLOATBUF0\[24\].A BYTE\[3\].FLOATBUF0\[24\].TE_B
+ VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG net236 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_60_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_110_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_83_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XA0BUF\[4\].__cell__ A0[4] VGND VGND VPWR VPWR A0BUF\[4\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV_123 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__inv_1
XFILLER_130_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XDIBUF\[32\].__cell__ Di0[32] VGND VGND VPWR VPWR DIBUF\[32\].X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_109_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_48_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_98_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_61_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_15_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_77_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CG net30 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_18_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_83_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_83_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV_155 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__inv_1
XFILLER_59_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_78_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG net143 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_128_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_53_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_130_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_124_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG net90 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_87_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[0\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_112_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[6\] Do0_REG.CLKBUF\[4\] BYTE\[4\].FLOATBUF0\[38\].Z
+ VGND VGND VPWR VPWR Do0[38] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG net247 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_26_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_21_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_1_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_76_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CLKINV_221 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__inv_1
XFILLER_84_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG net203 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_72_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_125_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_121_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_131_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_85_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_107_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_13_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CLKINV_125 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__inv_1
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_95_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDIBUF\[22\].__cell__ Di0[22] VGND VGND VPWR VPWR DIBUF\[22\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_51_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_112_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDIBUF\[61\].__cell__ Di0[61] VGND VGND VPWR VPWR DIBUF\[61\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[6\].FLOATBUF0\[49\].__cell__ BYTE\[6\].FLOATBUF0\[48\].A BYTE\[6\].FLOATBUF0\[48\].TE_B
+ VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_78_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_77_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_131_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[2\].FLOATBUF0\[17\].__cell__ BYTE\[2\].FLOATBUF0\[16\].A BYTE\[2\].FLOATBUF0\[16\].TE_B
+ VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG net101 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CLKINV_157 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__inv_1
XFILLER_48_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_24_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_32_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_101_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDIBUF\[6\].__cell__ Di0[6] VGND VGND VPWR VPWR DIBUF\[6\].X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_128_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_13_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG net214 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[5\].FLOATBUF0\[40\].__cell__ BYTE\[5\].FLOATBUF0\[40\].A BYTE\[5\].FLOATBUF0\[40\].TE_B
+ VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_14_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_13_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_68_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_83_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_124_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_120_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_74_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XWEBUF\[2\].__cell__ WE0[2] VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[2\].A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG net161 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_124_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[3\] Do0_REG.CLKBUF\[1\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VGND VGND VPWR VPWR Do0[11] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CG net8 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CLKINV_223 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_33_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV_250 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__inv_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_130_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_110_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV_1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__inv_1
XFILLER_56_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_61_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_133_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_7_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_116_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_97_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_103_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CLKINV_127 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__inv_1
XFILLER_102_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG net112 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_57_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_112_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_97_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_47_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG net68 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_63_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_62_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[12\].__cell__ Di0[12] VGND VGND VPWR VPWR DIBUF\[12\].X sky130_fd_sc_hd__clkbuf_16
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_125_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_97_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDIBUF\[51\].__cell__ Di0[51] VGND VGND VPWR VPWR DIBUF\[51\].X sky130_fd_sc_hd__clkbuf_16
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_26_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG net59 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_22_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_5_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_131_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV_129 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_17_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_83_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CLKINV_159 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__inv_1
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV_186 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_4_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_113_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG net172 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_112_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_37_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_73_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[3\] Do0_REG.CLKBUF\[6\] BYTE\[6\].FLOATBUF0\[51\].Z
+ VGND VGND VPWR VPWR Do0[51] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_89_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_94_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_60_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.DEC0.ABUF\[2\] A0BUF\[2\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.A_buf\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_41_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_126_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_63_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_73_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_108_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV_252 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__inv_1
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV_11 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__inv_1
XFILLER_92_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XDo0_REG.Do_CLKBUF\[5\] Do0_REG.CLK_buf VGND VGND VPWR VPWR Do0_REG.CLKBUF\[5\] sky130_fd_sc_hd__clkbuf_4
XFILLER_45_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_87_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XBYTE\[4\].FLOATBUF0\[32\].__cell__ BYTE\[4\].FLOATBUF0\[32\].A BYTE\[4\].FLOATBUF0\[32\].TE_B
+ VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG net79 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_105_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[7\] Do0_REG.CLKBUF\[2\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VGND VGND VPWR VPWR Do0[23] sky130_fd_sc_hd__dfxtp_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_7_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_78_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_77_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_65_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_61_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WEBUF\[0\].__cell__ SLICE\[0\].RAM8.WEBUF\[0\].A VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WEBUF\[0\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_119_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG net26 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_130_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XBYTE\[0\].FLOATBUF0\[5\].__cell__ BYTE\[0\].FLOATBUF0\[0\].A BYTE\[0\].FLOATBUF0\[0\].TE_B
+ VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG net183 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_120_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_90_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_128_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_109_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_3_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[41\].__cell__ Di0[41] VGND VGND VPWR VPWR DIBUF\[41\].X sky130_fd_sc_hd__clkbuf_16
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG net139 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WEBUF\[2\].__cell__ SLICE\[0\].RAM8.WEBUF\[2\].A VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WEBUF\[2\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV_188 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__inv_1
XFILLER_57_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_29_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CLKINV_29 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__inv_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_7_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_34_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[0\] Do0_REG.CLKBUF\[3\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VGND VGND VPWR VPWR Do0[24] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG net243 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_122_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_49_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WEBUF\[4\].__cell__ SLICE\[0\].RAM8.WEBUF\[4\].A VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WEBUF\[4\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_8_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_95_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_79_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_54_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CLKINV_254 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[7\] Do0_REG.CLKBUF\[7\] BYTE\[7\].FLOATBUF0\[63\].Z
+ VGND VGND VPWR VPWR Do0[63] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CG net37 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_104_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_89_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_18_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_40_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WEBUF\[6\].__cell__ SLICE\[0\].RAM8.WEBUF\[6\].A VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WEBUF\[6\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_24_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_59_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG net150 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_6_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_89_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_77_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_60_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[7\].FLOATBUF0\[56\].__cell__ BYTE\[7\].FLOATBUF0\[56\].A BYTE\[7\].FLOATBUF0\[56\].TE_B
+ VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_24_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[3\].FLOATBUF0\[24\].__cell__ BYTE\[3\].FLOATBUF0\[24\].A BYTE\[3\].FLOATBUF0\[24\].TE_B
+ VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG net97 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CLKINV_37 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_132_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV_49 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_70_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_42_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XA0BUF\[3\].__cell__ A0[3] VGND VGND VPWR VPWR A0BUF\[3\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_124_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG net254 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_124_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDIBUF\[31\].__cell__ Di0[31] VGND VGND VPWR VPWR DIBUF\[31\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_123_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_61_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_88_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG net210 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_84_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_44_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_90_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_128_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV_3 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_124_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CG net48 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_66_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_33_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_107_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CLKINV_141 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__inv_1
XFILLER_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG net4 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_72_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_72_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CLKINV_69 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__inv_1
XFILLER_133_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_121_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV_226 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__inv_1
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_70_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CLKINV_256 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__inv_1
XFILLER_7_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[4\] Do0_REG.CLKBUF\[4\] BYTE\[4\].FLOATBUF0\[36\].Z
+ VGND VGND VPWR VPWR Do0[36] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_53_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_88_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_131_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_29_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG net108 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_95_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_75_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_44_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_113_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.DEC0.AND0 SLICE\[2\].RAM8.DEC0.A_buf\[0\] SLICE\[2\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[0\].W.SEL0 sky130_fd_sc_hd__nor4b_2
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_66_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CLKINV_45 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__inv_1
XFILLER_34_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_108_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV_57 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__inv_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG net221 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_94_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_45_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_26_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_99_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_98_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_67_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_66_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_27_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CLKINV_111 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__inv_1
XFILLER_108_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[21\].__cell__ Di0[21] VGND VGND VPWR VPWR DIBUF\[21\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_108_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CG net15 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_92_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[60\].__cell__ Di0[60] VGND VGND VPWR VPWR DIBUF\[60\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_5_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_96_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XBYTE\[6\].FLOATBUF0\[48\].__cell__ BYTE\[6\].FLOATBUF0\[48\].A BYTE\[6\].FLOATBUF0\[48\].TE_B
+ VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XBYTE\[2\].FLOATBUF0\[16\].__cell__ BYTE\[2\].FLOATBUF0\[16\].A BYTE\[2\].FLOATBUF0\[16\].TE_B
+ VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_87_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CLKINV_77 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__inv_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV_89 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__inv_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_34_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_104_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_65_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CLKINV_143 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__inv_1
XFILLER_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV_170 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__inv_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG net119 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_114_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDIBUF\[5\].__cell__ Di0[5] VGND VGND VPWR VPWR DIBUF\[5\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_84_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTIE0\[7\].__cell__ VGND VGND VPWR VPWR TIE0\[7\].__cell__/HI BYTE\[7\].FLOATBUF0\[56\].A
+ sky130_fd_sc_hd__conb_1
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV_228 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG net75 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_106_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_120_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_74_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_74_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_112_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[1\] Do0_REG.CLKBUF\[1\] BYTE\[1\].FLOATBUF0\[9\].Z
+ VGND VGND VPWR VPWR Do0[9] sky130_fd_sc_hd__dfxtp_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG net232 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_66_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CLKINV_53 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__inv_1
XFILLER_111_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XWEBUF\[1\].__cell__ WE0[1] VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[1\].A sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_48_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_16_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG net179 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_131_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_98_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[7\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_34_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_57_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_17_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_53_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_9_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_107_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.DEC0.AND1 SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[0\] SLICE\[2\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[1\].W.SEL0 sky130_fd_sc_hd__and4bb_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_108_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_118_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[11\].__cell__ Di0[11] VGND VGND VPWR VPWR DIBUF\[11\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_123_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CLKINV_85 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__inv_1
XFILLER_103_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV_97 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__inv_1
XFILLER_13_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDIBUF\[50\].__cell__ Di0[50] VGND VGND VPWR VPWR DIBUF\[50\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_126_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG net86 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_110_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_63_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_6_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV_172 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__inv_1
XFILLER_2_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_104_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[1\] Do0_REG.CLKBUF\[6\] BYTE\[6\].FLOATBUF0\[49\].Z
+ VGND VGND VPWR VPWR Do0[49] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_73_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG net199 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG net33 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.DEC0.ABUF\[0\] A0BUF\[0\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.A_buf\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_96_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG net190 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CLKINV_61 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_117_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG net146 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_109_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_93_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.Do_CLKBUF\[3\] Do0_REG.CLK_buf VGND VGND VPWR VPWR Do0_REG.CLKBUF\[3\] sky130_fd_sc_hd__clkbuf_4
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_96_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_96_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFBUFENBUF0\[7\].__cell__ EN0 VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].TE_B sky130_fd_sc_hd__clkbuf_2
XFILLER_71_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_75_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_101_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_47_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[5\] Do0_REG.CLKBUF\[2\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VGND VGND VPWR VPWR Do0[21] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_55_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_124_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[6\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG net250 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CLKINV_5 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CLKINV_93 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__inv_1
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_121_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_47_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_112_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[0\].FLOATBUF0\[4\].__cell__ BYTE\[0\].FLOATBUF0\[0\].A BYTE\[0\].FLOATBUF0\[0\].TE_B
+ VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_22_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG net44 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_30_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_116_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_89_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_72_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[40\].__cell__ Di0[40] VGND VGND VPWR VPWR DIBUF\[40\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_35_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WEBUF\[1\].__cell__ SLICE\[0\].RAM8.WEBUF\[1\].A VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WEBUF\[1\].X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_31_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_129_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG net157 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_7_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_98_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.DEC0.AND2 SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[1\] SLICE\[2\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[2\].W.SEL0 sky130_fd_sc_hd__and4bb_2
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CLKINV_174 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__inv_1
XFILLER_93_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_123_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_116_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_104_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_84_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_9_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_105_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WEBUF\[3\].__cell__ SLICE\[0\].RAM8.WEBUF\[3\].A VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WEBUF\[3\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_99_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[5\] Do0_REG.CLKBUF\[7\] BYTE\[7\].FLOATBUF0\[61\].Z
+ VGND VGND VPWR VPWR Do0[61] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_23_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_92_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_57_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_9_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG net217 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_107_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV_210 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_76_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CLKINV_240 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__inv_1
XFILLER_63_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_55_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CG net55 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WEBUF\[5\].__cell__ SLICE\[0\].RAM8.WEBUF\[5\].A VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WEBUF\[5\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[5\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_61_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG net11 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.DEC0.ABUF\[1\] A0BUF\[1\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.A_buf\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_115_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV_114 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__inv_1
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_106_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG net168 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_114_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_120_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_87_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_115_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_96_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XA0BUF\[2\].__cell__ A0[2] VGND VGND VPWR VPWR A0BUF\[2\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG net115 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDIBUF\[30\].__cell__ Di0[30] VGND VGND VPWR VPWR DIBUF\[30\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_80_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV_146 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__inv_1
XFILLER_75_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_75_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CLKINV_176 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__inv_1
XFILLER_71_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_31_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_93_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG net228 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_131_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_83_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_107_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_121_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC0.AND3 SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[0\] SLICE\[2\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[3\].W.SEL0 sky130_fd_sc_hd__and4b_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[2\] Do0_REG.CLKBUF\[4\] BYTE\[4\].FLOATBUF0\[34\].Z
+ VGND VGND VPWR VPWR Do0[34] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CG net22 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_118_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV_212 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_41_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_43_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_68_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_75_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_91_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_31_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_113_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG net135 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_123_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_89_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_100_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[4\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG net126 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV_116 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__inv_1
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_122_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_24_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG net82 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[6\] Do0_REG.CLKBUF\[0\] BYTE\[0\].FLOATBUF0\[6\].Z
+ VGND VGND VPWR VPWR Do0[6] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_86_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_10_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG net239 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_108_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_2_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_33_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_60_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_81_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_114_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG net195 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_68_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_64_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV_148 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__inv_1
XDIBUF\[20\].__cell__ Di0[20] VGND VGND VPWR VPWR DIBUF\[20\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_101_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG net186 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_124_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_93_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_119_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_4_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDIBUF\[4\].__cell__ Di0[4] VGND VGND VPWR VPWR DIBUF\[4\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTIE0\[6\].__cell__ VGND VGND VPWR VPWR TIE0\[6\].__cell__/HI BYTE\[6\].FLOATBUF0\[48\].A
+ sky130_fd_sc_hd__conb_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_124_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CLKINV_7 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__inv_1
XFILLER_53_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_46_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CLKINV_214 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__inv_1
XFILLER_128_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV_241 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__inv_1
XFILLER_69_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG net93 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_32_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.DEC0.ENBUF SLICE\[1\].RAM8.DEC0.EN VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.EN_buf
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_63_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_73_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_43_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_129_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[6\] Do0_REG.CLKBUF\[5\] BYTE\[5\].FLOATBUF0\[46\].Z
+ VGND VGND VPWR VPWR Do0[46] sky130_fd_sc_hd__dfxtp_1
XWEBUF\[0\].__cell__ WE0[0] VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[0\].A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_112_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.DEC0.AND4 SLICE\[2\].RAM8.DEC0.A_buf\[0\] SLICE\[2\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[4\].W.SEL0 sky130_fd_sc_hd__and4bb_2
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_94_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG net206 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_104_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CLKINV_118 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__inv_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[3\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_25_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_76_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_90_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_98_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_58_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_67_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV_10 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__inv_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG net153 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_89_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_92_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_122_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV_177 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_83_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_64_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[10\].__cell__ Di0[10] VGND VGND VPWR VPWR DIBUF\[10\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_32_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_87_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_131_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_11_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_10_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_124_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_65_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG net104 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_127_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_83_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_64_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_42_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CLKINV_16 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CLKINV_216 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__inv_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG net51 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_120_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV_28 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV_243 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__inv_1
XFILLER_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.Do_CLKBUF\[1\] Do0_REG.CLK_buf VGND VGND VPWR VPWR Do0_REG.CLKBUF\[1\] sky130_fd_sc_hd__clkbuf_4
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_61_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_14_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_128_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_111_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_25_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[3\] Do0_REG.CLKBUF\[2\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VGND VGND VPWR VPWR Do0[19] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG net164 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_43_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFBUFENBUF0\[6\].__cell__ EN0 VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].TE_B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_7_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_131_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_130_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[2\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_72_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_13_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_75_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.DEC0.AND5 SLICE\[2\].RAM8.DEC0.A_buf\[1\] SLICE\[2\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[5\].W.SEL0 sky130_fd_sc_hd__and4b_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_47_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.DEC0.ABUF\[2\] A0BUF\[2\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.A_buf\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_50_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV_179 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__inv_1
XFILLER_72_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_26_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_41_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_40_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XBYTE\[0\].FLOATBUF0\[3\].__cell__ BYTE\[0\].FLOATBUF0\[0\].A BYTE\[0\].FLOATBUF0\[0\].TE_B
+ VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG net71 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_110_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_88_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_124_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_86_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CG net62 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_129_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_116_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WEBUF\[0\].__cell__ SLICE\[0\].RAM8.WEBUF\[0\].A VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WEBUF\[0\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_18_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG net18 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_45_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CLKINV_24 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__inv_1
XFILLER_41_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.Root_CLKBUF CLKBUF.X VGND VGND VPWR VPWR Do0_REG.CLK_buf sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV_130 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__inv_1
XFILLER_5_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV_36 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__inv_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_96_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_110_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CLKINV_160 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_95_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_44_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG net175 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_20_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_101_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[3\] Do0_REG.CLKBUF\[7\] BYTE\[7\].FLOATBUF0\[59\].Z
+ VGND VGND VPWR VPWR Do0[59] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_23_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CLKINV_245 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG net131 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_123_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WEBUF\[2\].__cell__ SLICE\[0\].RAM8.WEBUF\[2\].A VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WEBUF\[2\].X sky130_fd_sc_hd__clkbuf_2
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_127_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG net122 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_51_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_2_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_65_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_92_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG net235 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_41_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV_68 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WEBUF\[4\].__cell__ SLICE\[0\].RAM8.WEBUF\[4\].A VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WEBUF\[4\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[1\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_84_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[7\] Do0_REG.CLKBUF\[3\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VGND VGND VPWR VPWR Do0[31] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_114_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_3_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_3_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_87_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.genblk1.CG net29 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV_100 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__inv_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_53_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_80_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_40_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_122_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CLKINV_32 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__inv_1
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV_44 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__inv_1
XFILLER_8_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XA0BUF\[1\].__cell__ A0[1] VGND VGND VPWR VPWR A0BUF\[1\].X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG net142 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_125_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.DEC0.AND6 SLICE\[2\].RAM8.DEC0.A_buf\[0\] SLICE\[2\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[6\].W.SEL0 sky130_fd_sc_hd__and4b_2
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_35_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_104_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_116_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_103_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV_132 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__inv_1
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_13_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG net89 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_91_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_44_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_32_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV_217 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__inv_1
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CLKINV_247 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__inv_1
XFILLER_99_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[0\] Do0_REG.CLKBUF\[4\] BYTE\[4\].FLOATBUF0\[32\].Z
+ VGND VGND VPWR VPWR Do0[32] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG net246 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_104_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_57_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_85_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG net202 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_13_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_127_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_5_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV_76 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_118_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_86_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_55_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_27_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CG net40 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_35_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_40_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_121_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_123_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[0\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_92_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_91_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_91_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[4\] Do0_REG.CLKBUF\[0\] BYTE\[0\].FLOATBUF0\[4\].Z
+ VGND VGND VPWR VPWR Do0[4] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_87_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_101_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_87_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_101_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_129_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CLKINV_40 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__inv_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CLKINV_102 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__inv_1
XFILLER_3_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_3_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV_52 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__inv_1
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_130_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG net100 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_40_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_121_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_102_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_46_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_70_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_109_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_81_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CLKINV_134 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG net213 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV_161 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__inv_1
XFILLER_116_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CLKINV_191 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV_219 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__inv_1
XFILLER_106_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_102_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_78_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CLKINV_72 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_98_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV_84 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__inv_1
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.DEC0.AND7 SLICE\[2\].RAM8.DEC0.A_buf\[0\] SLICE\[2\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WORD\[7\].W.SEL0 sky130_fd_sc_hd__and4_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_54_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.DEC0.AND0 SLICE\[0\].RAM8.DEC0.A_buf\[0\] SLICE\[0\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[0\].W.SEL0 sky130_fd_sc_hd__nor4b_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CG net7 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_30_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[3\].__cell__ Di0[3] VGND VGND VPWR VPWR DIBUF\[3\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_85_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_26_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTIE0\[5\].__cell__ VGND VGND VPWR VPWR TIE0\[5\].__cell__/HI BYTE\[5\].FLOATBUF0\[40\].A
+ sky130_fd_sc_hd__conb_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV_193 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__inv_1
XFILLER_41_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_40_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_129_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[4\] Do0_REG.CLKBUF\[5\] BYTE\[5\].FLOATBUF0\[44\].Z
+ VGND VGND VPWR VPWR Do0[44] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CLKINV_200 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__inv_1
XFILLER_99_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_125_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_90_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_10_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_116_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG net111 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV_60 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_88_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG net67 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_72_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_71_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.genblk1.CLKINV_104 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_67_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG net224 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_109_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG net58 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_46_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_60_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_84_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_36_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG net171 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_59_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CLKINV_136 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_104_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[7\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV_163 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__inv_1
XFILLER_59_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDIBUF\[59\].__cell__ Di0[59] VGND VGND VPWR VPWR DIBUF\[59\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_74_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CLKINV_80 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__inv_1
XFILLER_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV_92 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_127_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_110_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_108_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_71_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_43_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_124_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV_195 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__inv_1
XFILLER_30_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_130_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_40_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG net78 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_107_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_121_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_87_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[1\] Do0_REG.CLKBUF\[2\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VGND VGND VPWR VPWR Do0[17] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_44_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_125_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_79_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_19_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.DEC0.AND1 SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[0\] SLICE\[0\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[1\].W.SEL0 sky130_fd_sc_hd__and4bb_2
XFILLER_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_104_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG net25 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_85_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFBUFENBUF0\[5\].__cell__ EN0 VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].TE_B sky130_fd_sc_hd__clkbuf_2
XFILLER_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_68_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_76_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG net182 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_48_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_76_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_117_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_99_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG net138 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.DEC0.ABUF\[0\] A0BUF\[0\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.A_buf\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_129_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_116_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_104_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_95_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XBYTE\[7\].FLOATBUF0\[63\].__cell__ BYTE\[7\].FLOATBUF0\[56\].A BYTE\[7\].FLOATBUF0\[56\].TE_B
+ VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_49_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_99_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XBYTE\[3\].FLOATBUF0\[31\].__cell__ BYTE\[3\].FLOATBUF0\[24\].A BYTE\[3\].FLOATBUF0\[24\].TE_B
+ VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XBYTE\[0\].FLOATBUF0\[2\].__cell__ BYTE\[0\].FLOATBUF0\[0\].A BYTE\[0\].FLOATBUF0\[0\].TE_B
+ VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CLKINV_165 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__inv_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_104_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[6\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG net242 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_132_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_105_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[49\].__cell__ Di0[49] VGND VGND VPWR VPWR DIBUF\[49\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_121_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_5_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_123_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_110_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[1\] Do0_REG.CLKBUF\[7\] BYTE\[7\].FLOATBUF0\[57\].Z
+ VGND VGND VPWR VPWR Do0[57] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_51_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_3_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_105_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG net36 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_78_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CLKINV_197 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__inv_1
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_76_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_111_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_69_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_65_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_37_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV_201 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__inv_1
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CLKINV_231 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_99_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WEBUF\[1\].__cell__ SLICE\[0\].RAM8.WEBUF\[1\].A VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WEBUF\[1\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG net149 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_71_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_74_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_61_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_15_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_30_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_116_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_97_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.CLKBUF.__cell__ CLKBUF.X VGND VGND VPWR VPWR SLICE\[3\].RAM8.CLKBUF.X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_52_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV_105 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__inv_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_107_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[5\] Do0_REG.CLKBUF\[3\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VGND VGND VPWR VPWR Do0[29] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_121_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_29_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_113_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_44_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WEBUF\[3\].__cell__ SLICE\[0\].RAM8.WEBUF\[3\].A VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WEBUF\[3\].X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_12_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_12_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_121_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG net253 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_93_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.DEC0.AND2 SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[1\] SLICE\[0\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[2\].W.SEL0 sky130_fd_sc_hd__and4bb_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_34_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_85_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG net209 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_26_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_103_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV_137 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__inv_1
XFILLER_71_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CLKINV_167 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_8_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_125_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_67_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CG net47 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_31_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[5\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_116_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDIBUF\[39\].__cell__ Di0[39] VGND VGND VPWR VPWR DIBUF\[39\].X sky130_fd_sc_hd__clkbuf_16
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG net3 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XA0BUF\[0\].__cell__ A0[0] VGND VGND VPWR VPWR A0BUF\[0\].X sky130_fd_sc_hd__clkbuf_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_110_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG net160 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_9_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XBYTE\[6\].FLOATBUF0\[55\].__cell__ BYTE\[6\].FLOATBUF0\[48\].A BYTE\[6\].FLOATBUF0\[48\].TE_B
+ VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_132_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_82_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CLKINV_199 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__inv_1
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XBYTE\[2\].FLOATBUF0\[23\].__cell__ BYTE\[2\].FLOATBUF0\[16\].A BYTE\[2\].FLOATBUF0\[16\].TE_B
+ VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV_203 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__inv_1
XFILLER_127_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG net107 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_6_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_9_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_114_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG net220 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_92_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV_107 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_2_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[2\] Do0_REG.CLKBUF\[0\] BYTE\[0\].FLOATBUF0\[2\].Z
+ VGND VGND VPWR VPWR Do0[2] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_119_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_87_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_75_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_109_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_127_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_46_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CG net14 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XCLKBUF.__cell__ CLK VGND VGND VPWR VPWR CLKBUF.X sky130_fd_sc_hd__clkbuf_4
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_96_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_96_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_84_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_53_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV_139 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV_19 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__inv_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_121_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_12_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_8_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_81_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.DEC0.AND3 SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[0\] SLICE\[0\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[3\].W.SEL0 sky130_fd_sc_hd__and4b_2
XFILLER_22_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_42_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[4\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG net118 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XDIBUF\[29\].__cell__ Di0[29] VGND VGND VPWR VPWR DIBUF\[29\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_112_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_13_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_107_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_68_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.CLKBUF.__cell__ CLKBUF.X VGND VGND VPWR VPWR SLICE\[1\].RAM8.CLKBUF.X
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG net74 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_84_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_67_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG net231 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_81_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CLKINV_205 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__inv_1
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_73_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_5_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_122_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_49_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_32_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XDIBUF\[2\].__cell__ Di0[2] VGND VGND VPWR VPWR DIBUF\[2\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_12_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[2\] Do0_REG.CLKBUF\[5\] BYTE\[5\].FLOATBUF0\[42\].Z
+ VGND VGND VPWR VPWR Do0[42] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG net178 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTIE0\[4\].__cell__ VGND VGND VPWR VPWR TIE0\[4\].__cell__/HI BYTE\[4\].FLOATBUF0\[32\].A
+ sky130_fd_sc_hd__conb_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_99_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[5\].FLOATBUF0\[47\].__cell__ BYTE\[5\].FLOATBUF0\[40\].A BYTE\[5\].FLOATBUF0\[40\].TE_B
+ VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_82_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[1\].FLOATBUF0\[15\].__cell__ BYTE\[1\].FLOATBUF0\[10\].A BYTE\[1\].FLOATBUF0\[10\].TE_B
+ VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CLKINV_109 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__inv_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_10_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_110_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_76_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CLKINV_15 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_67_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV_27 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_23_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_3_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_76_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_10_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[6\] Do0_REG.CLKBUF\[1\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VGND VGND VPWR VPWR Do0[14] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG net85 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_60_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_20_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_102_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_11_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_11_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_87_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_120_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_47_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_62_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG net198 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[1\].FLOATBUF0\[9\].__cell__ BYTE\[1\].FLOATBUF0\[10\].A BYTE\[1\].FLOATBUF0\[10\].TE_B
+ VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[3\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[19\].__cell__ Di0[19] VGND VGND VPWR VPWR DIBUF\[19\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_69_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_65_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[58\].__cell__ Di0[58] VGND VGND VPWR VPWR DIBUF\[58\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_106_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG net189 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_102_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_98_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG net145 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_121_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CLKINV_207 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__inv_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.DEC0.AND4 SLICE\[0\].RAM8.DEC0.A_buf\[0\] SLICE\[0\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[4\].W.SEL0 sky130_fd_sc_hd__and4bb_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV_234 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__inv_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_116_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_84_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_34_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_107_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_35_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CLKINV_23 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG net249 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_131_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV_35 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG net96 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_26_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_110_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_5_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[6\] Do0_REG.CLKBUF\[6\] BYTE\[6\].FLOATBUF0\[54\].Z
+ VGND VGND VPWR VPWR Do0[54] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_48_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_95_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_13_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFBUFENBUF0\[4\].__cell__ EN0 VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].TE_B sky130_fd_sc_hd__clkbuf_2
XFILLER_117_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG net43 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XBYTE\[4\].FLOATBUF0\[39\].__cell__ BYTE\[4\].FLOATBUF0\[32\].A BYTE\[4\].FLOATBUF0\[32\].TE_B
+ VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_131_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_100_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_107_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG net156 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_113_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WEBUF\[7\].__cell__ SLICE\[0\].RAM8.WEBUF\[7\].A VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WEBUF\[7\].X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_82_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[7\].FLOATBUF0\[62\].__cell__ BYTE\[7\].FLOATBUF0\[56\].A BYTE\[7\].FLOATBUF0\[56\].TE_B
+ VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_104_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_132_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV_67 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_59_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_86_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_46_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_14_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBYTE\[3\].FLOATBUF0\[30\].__cell__ BYTE\[3\].FLOATBUF0\[24\].A BYTE\[3\].FLOATBUF0\[24\].TE_B
+ VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z sky130_fd_sc_hd__ebufn_2
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[2\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[0\].FLOATBUF0\[1\].__cell__ BYTE\[0\].FLOATBUF0\[0\].A BYTE\[0\].FLOATBUF0\[0\].TE_B
+ VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_110_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CLKINV_151 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDIBUF\[48\].__cell__ Di0[48] VGND VGND VPWR VPWR DIBUF\[48\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_24_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV_236 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__inv_1
XFILLER_118_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CLKINV_31 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__inv_1
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV_43 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__inv_1
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_83_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_12_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.DEC0.ABUF\[2\] A0BUF\[2\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.A_buf\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_8_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CG net54 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_125_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_121_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_94_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_47_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WEBUF\[0\].__cell__ SLICE\[0\].RAM8.WEBUF\[0\].A VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WEBUF\[0\].X sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.DEC0.AND5 SLICE\[0\].RAM8.DEC0.A_buf\[1\] SLICE\[0\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[5\].W.SEL0 sky130_fd_sc_hd__and4b_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_128_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG net10 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_53_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_119_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[3\] Do0_REG.CLKBUF\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VGND VGND VPWR VPWR Do0[27] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_108_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG net167 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_104_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WEBUF\[2\].__cell__ SLICE\[0\].RAM8.WEBUF\[2\].A VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WEBUF\[2\].X sky130_fd_sc_hd__clkbuf_2
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG net114 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_22_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV_75 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__inv_1
XFILLER_21_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_5_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_79_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_103_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_72_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_44_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_94_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_50_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_117_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG net227 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_22_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[1\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV_180 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__inv_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_77_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_72_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_9_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[38\].__cell__ Di0[38] VGND VGND VPWR VPWR DIBUF\[38\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_5_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_113_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CLKINV_238 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV_51 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__inv_1
XFILLER_28_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CG net21 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_105_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_100_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[6\].FLOATBUF0\[54\].__cell__ BYTE\[6\].FLOATBUF0\[48\].A BYTE\[6\].FLOATBUF0\[48\].TE_B
+ VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_2_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[2\].FLOATBUF0\[22\].__cell__ BYTE\[2\].FLOATBUF0\[16\].A BYTE\[2\].FLOATBUF0\[16\].TE_B
+ VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG net134 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_102_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_78_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG net125 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_128_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_123_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_111_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[0\] Do0_REG.CLKBUF\[0\] BYTE\[0\].FLOATBUF0\[0\].Z
+ VGND VGND VPWR VPWR Do0[0] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG net81 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_107_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.genblk1.CLKINV_71 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV_83 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG net238 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_120_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDEC0.AND0 A0BUF\[3\].X A0BUF\[4\].X DEC0.EN VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.EN
+ sky130_fd_sc_hd__nor3b_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.DEC0.AND6 SLICE\[0\].RAM8.DEC0.A_buf\[0\] SLICE\[0\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[6\].W.SEL0 sky130_fd_sc_hd__and4b_2
XFILLER_15_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_128_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG net194 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[7\] Do0_REG.CLKBUF\[4\] BYTE\[4\].FLOATBUF0\[39\].Z
+ VGND VGND VPWR VPWR Do0[39] sky130_fd_sc_hd__dfxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_102_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG net185 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CG net32 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_79_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_94_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_43_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_116_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_112_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_65_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CLKINV_182 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__inv_1
XFILLER_26_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_80_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[0\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_107_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_115_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_17_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[28\].__cell__ Di0[28] VGND VGND VPWR VPWR DIBUF\[28\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_79_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_117_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_85_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG net92 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_123_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_29_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[0\] Do0_REG.CLKBUF\[5\] BYTE\[5\].FLOATBUF0\[40\].Z
+ VGND VGND VPWR VPWR Do0[40] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV_91 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__inv_1
XFILLER_117_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_105_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[1\].__cell__ Di0[1] VGND VGND VPWR VPWR DIBUF\[1\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG net205 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_100_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_86_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XTIE0\[3\].__cell__ VGND VGND VPWR VPWR TIE0\[3\].__cell__/HI BYTE\[3\].FLOATBUF0\[24\].A
+ sky130_fd_sc_hd__conb_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_22_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_128_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[5\].FLOATBUF0\[46\].__cell__ BYTE\[5\].FLOATBUF0\[40\].A BYTE\[5\].FLOATBUF0\[40\].TE_B
+ VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_2_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV_9 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__inv_1
XFILLER_111_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_77_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[1\].FLOATBUF0\[14\].__cell__ BYTE\[1\].FLOATBUF0\[10\].A BYTE\[1\].FLOATBUF0\[10\].TE_B
+ VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_110_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV_122 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_59_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_128_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[4\] Do0_REG.CLKBUF\[1\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VGND VGND VPWR VPWR Do0[12] sky130_fd_sc_hd__dfxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_123_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_46_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_119_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_106_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV_154 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__inv_1
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XDEC0.AND1 A0BUF\[4\].X A0BUF\[3\].X DEC0.EN VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.EN
+ sky130_fd_sc_hd__and3b_2
XFILLER_28_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.DEC0.AND7 SLICE\[0\].RAM8.DEC0.A_buf\[0\] SLICE\[0\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WORD\[7\].W.SEL0 sky130_fd_sc_hd__and4_2
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CLKINV_184 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__inv_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG net103 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_97_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_108_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XBYTE\[1\].FLOATBUF0\[8\].__cell__ BYTE\[1\].FLOATBUF0\[10\].A BYTE\[1\].FLOATBUF0\[10\].TE_B
+ VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[18\].__cell__ Di0[18] VGND VGND VPWR VPWR DIBUF\[18\].X sky130_fd_sc_hd__clkbuf_16
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_121_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[57\].__cell__ Di0[57] VGND VGND VPWR VPWR DIBUF\[57\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG net216 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_58_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG net50 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_47_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_122_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_89_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_130_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_57_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV_220 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG net163 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_8_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_60_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_95_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[7\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_86_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_81_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_14_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_10_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_122_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[4\] Do0_REG.CLKBUF\[6\] BYTE\[6\].FLOATBUF0\[52\].Z
+ VGND VGND VPWR VPWR Do0[52] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_60_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.DEC0.AND0 SLICE\[3\].RAM8.DEC0.A_buf\[0\] SLICE\[3\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[0\].W.SEL0 sky130_fd_sc_hd__nor4b_2
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_9_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV_124 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__inv_1
XFILLER_114_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_68_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_51_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_90_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_132_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFBUFENBUF0\[3\].__cell__ EN0 VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].TE_B sky130_fd_sc_hd__clkbuf_2
XFILLER_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_128_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_123_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG net70 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_2_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XBYTE\[4\].FLOATBUF0\[38\].__cell__ BYTE\[4\].FLOATBUF0\[32\].A BYTE\[4\].FLOATBUF0\[32\].TE_B
+ VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.Do_CLKBUF\[6\] Do0_REG.CLK_buf VGND VGND VPWR VPWR Do0_REG.CLKBUF\[6\] sky130_fd_sc_hd__clkbuf_4
XFILLER_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_127_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_87_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_102_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CG net61 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV_156 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__inv_1
XFILLER_109_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_3_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_105_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_132_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG net17 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WEBUF\[6\].__cell__ SLICE\[0\].RAM8.WEBUF\[6\].A VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WEBUF\[6\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_108_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_69_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XBYTE\[7\].FLOATBUF0\[61\].__cell__ BYTE\[7\].FLOATBUF0\[56\].A BYTE\[7\].FLOATBUF0\[56\].TE_B
+ VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_53_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG net174 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_9_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_68_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[0\].FLOATBUF0\[0\].__cell__ BYTE\[0\].FLOATBUF0\[0\].A BYTE\[0\].FLOATBUF0\[0\].TE_B
+ VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_24_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_98_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG net130 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_120_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[47\].__cell__ Di0[47] VGND VGND VPWR VPWR DIBUF\[47\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_101_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC0.AND2 A0BUF\[3\].X A0BUF\[4\].X DEC0.EN VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.EN
+ sky130_fd_sc_hd__and3b_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_128_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_97_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG net121 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_93_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_53_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CLKINV_222 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_44_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.DEC0.ABUF\[0\] A0BUF\[0\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.DEC0.A_buf\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_75_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[6\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_15_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG net234 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_110_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_119_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[1\] Do0_REG.CLKBUF\[3\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VGND VGND VPWR VPWR Do0[25] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_91_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CLKINV_126 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__inv_1
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_13_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_12_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_121_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG net28 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_129_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_85_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_76_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_91_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_57_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WEBUF\[1\].__cell__ SLICE\[0\].RAM8.WEBUF\[1\].A VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WEBUF\[1\].X sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.DEC0.AND1 SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[0\] SLICE\[3\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[1\].W.SEL0 sky130_fd_sc_hd__and4bb_2
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CLKINV_158 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__inv_1
XFILLER_5_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG net141 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_95_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_68_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV_185 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__inv_1
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_116_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_54_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_123_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_92_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_114_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_110_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_110_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG net245 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_118_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_3_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XDIBUF\[37\].__cell__ Di0[37] VGND VGND VPWR VPWR DIBUF\[37\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_19_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_15_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG net201 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_6_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_108_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV_18 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CLKINV_224 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__inv_1
XFILLER_37_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV_251 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[6\].FLOATBUF0\[53\].__cell__ BYTE\[6\].FLOATBUF0\[48\].A BYTE\[6\].FLOATBUF0\[48\].TE_B
+ VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_114_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_96_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[2\].FLOATBUF0\[21\].__cell__ BYTE\[2\].FLOATBUF0\[16\].A BYTE\[2\].FLOATBUF0\[16\].TE_B
+ VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CG net39 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_11_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.AND3 A0BUF\[4\].X A0BUF\[3\].X DEC0.EN VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.EN
+ sky130_fd_sc_hd__and3_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[5\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_10_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_124_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_97_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_18_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CLKINV_128 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__inv_1
XFILLER_21_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_107_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG net152 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_103_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_40_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_74_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[5\] Do0_REG.CLKBUF\[4\] BYTE\[4\].FLOATBUF0\[37\].Z
+ VGND VGND VPWR VPWR Do0[37] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_66_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG net99 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_22_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_89_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_103_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_57_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV_187 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__inv_1
XFILLER_13_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_13_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG net256 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG net212 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_100_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_34_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_108_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_122_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CLKINV_14 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV_26 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__inv_1
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.DEC0.AND2 SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[1\] SLICE\[3\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[2\].W.SEL0 sky130_fd_sc_hd__and4bb_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_121_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_50_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV_2 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CG net6 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDIBUF\[27\].__cell__ Di0[27] VGND VGND VPWR VPWR DIBUF\[27\].X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_74_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_6_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CLKINV_253 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__inv_1
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_77_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_95_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_64_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_48_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_24_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_132_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[4\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG net110 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_10_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_123_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_92_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_61_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG net66 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_60_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[0\].__cell__ Di0[0] VGND VGND VPWR VPWR DIBUF\[0\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_127_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XTIE0\[2\].__cell__ VGND VGND VPWR VPWR TIE0\[2\].__cell__/HI BYTE\[2\].FLOATBUF0\[16\].A
+ sky130_fd_sc_hd__conb_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XBYTE\[5\].FLOATBUF0\[45\].__cell__ BYTE\[5\].FLOATBUF0\[40\].A BYTE\[5\].FLOATBUF0\[40\].TE_B
+ VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_24_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG net223 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG net57 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_133_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[1\].FLOATBUF0\[13\].__cell__ BYTE\[1\].FLOATBUF0\[10\].A BYTE\[1\].FLOATBUF0\[10\].TE_B
+ VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_87_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_19_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[2\] Do0_REG.CLKBUF\[1\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VGND VGND VPWR VPWR Do0[10] sky130_fd_sc_hd__dfxtp_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_120_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XWEBUF\[7\].__cell__ WE0[7] VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[7\].A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.genblk1.CLKINV_189 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__inv_1
XFILLER_130_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG net170 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.genblk1.CLKINV_22 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__inv_1
XFILLER_33_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_116_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_106_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV_34 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_102_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_116_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_112_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_53_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_119_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_69_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV_140 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_44_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_109_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_121_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV_225 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__inv_1
XFILLER_116_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDIBUF\[17\].__cell__ Di0[17] VGND VGND VPWR VPWR DIBUF\[17\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_112_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.genblk1.CLKINV_255 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__inv_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG net77 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_10_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDIBUF\[56\].__cell__ Di0[56] VGND VGND VPWR VPWR DIBUF\[56\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_108_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_49_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.DEC0.AND3 SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[0\] SLICE\[3\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[3\].W.SEL0 sky130_fd_sc_hd__and4b_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV_66 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__inv_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_48_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_104_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_58_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[3\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_39_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[2\] Do0_REG.CLKBUF\[6\] BYTE\[6\].FLOATBUF0\[50\].Z
+ VGND VGND VPWR VPWR Do0[50] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.DEC0.ENBUF SLICE\[2\].RAM8.DEC0.EN VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.EN_buf
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_65_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG net181 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.DEC0.ABUF\[1\] A0BUF\[1\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.DEC0.A_buf\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_127_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_49_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG net137 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.genblk1.CLKINV_30 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__inv_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_128_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV_42 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__inv_1
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CLKINV_110 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__inv_1
XFILLER_117_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.Do_CLKBUF\[4\] Do0_REG.CLK_buf VGND VGND VPWR VPWR Do0_REG.CLKBUF\[4\] sky130_fd_sc_hd__clkbuf_4
XFILLER_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFBUFENBUF0\[2\].__cell__ EN0 VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].TE_B sky130_fd_sc_hd__clkbuf_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_114_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_130_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_110_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_56_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_71_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XBYTE\[4\].FLOATBUF0\[37\].__cell__ BYTE\[4\].FLOATBUF0\[32\].A BYTE\[4\].FLOATBUF0\[32\].TE_B
+ VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_47_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG net241 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_27_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[6\] Do0_REG.CLKBUF\[2\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VGND VGND VPWR VPWR Do0[22] sky130_fd_sc_hd__dfxtp_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_70_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG net88 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_7_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_73_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.genblk1.CLKINV_142 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_88_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WEBUF\[5\].__cell__ SLICE\[0\].RAM8.WEBUF\[5\].A VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WEBUF\[5\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XBYTE\[7\].FLOATBUF0\[60\].__cell__ BYTE\[7\].FLOATBUF0\[56\].A BYTE\[7\].FLOATBUF0\[56\].TE_B
+ VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_20_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV_227 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_87_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG net35 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_114_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV_74 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__inv_1
XFILLER_30_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CLKINV_48 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG net192 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XDIBUF\[46\].__cell__ Di0[46] VGND VGND VPWR VPWR DIBUF\[46\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_88_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_89_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[55\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_37_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_13_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WEBUF\[7\].__cell__ SLICE\[0\].RAM8.WEBUF\[7\].A VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WEBUF\[7\].X sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG net148 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_100_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_67_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_54_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[2\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_89_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_57_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV_50 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__inv_1
XFILLER_55_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.DEC0.AND4 SLICE\[3\].RAM8.DEC0.A_buf\[0\] SLICE\[3\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[4\].W.SEL0 sky130_fd_sc_hd__and4bb_2
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_96_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_67_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG net252 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_83_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_36_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_59_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_100_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.genblk1.CLKINV_112 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__inv_1
XFILLER_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[6\] Do0_REG.CLKBUF\[7\] BYTE\[7\].FLOATBUF0\[62\].Z
+ VGND VGND VPWR VPWR Do0[62] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_2_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[3\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_49_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV_4 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__inv_1
XFILLER_64_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_127_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_68_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.genblk1.CG net46 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_64_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_127_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WEBUF\[0\].__cell__ SLICE\[0\].RAM8.WEBUF\[0\].A VGND VGND VPWR VPWR
+ SLICE\[0\].RAM8.WEBUF\[0\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_98_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG net2 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_108_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_109_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CLKINV_70 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CLKINV_144 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__inv_1
XFILLER_123_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_77_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV_171 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__inv_1
XFILLER_92_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV_82 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_46_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_93_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG net159 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_119_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.DEC0.ABUF\[2\] A0BUF\[2\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.A_buf\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_127_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CLKINV_56 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CLKINV_229 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__inv_1
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_52_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_20_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XBYTE\[3\].FLOATBUF0\[29\].__cell__ BYTE\[3\].FLOATBUF0\[24\].A BYTE\[3\].FLOATBUF0\[24\].TE_B
+ VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_70_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_30_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG net106 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_34_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDIBUF\[36\].__cell__ Di0[36] VGND VGND VPWR VPWR DIBUF\[36\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_14_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_115_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_130_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_68_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_121_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_75_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[6\].FLOATBUF0\[52\].__cell__ BYTE\[6\].FLOATBUF0\[48\].A BYTE\[6\].FLOATBUF0\[48\].TE_B
+ VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_58_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_74_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG net219 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_124_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[2\].FLOATBUF0\[20\].__cell__ BYTE\[2\].FLOATBUF0\[16\].A BYTE\[2\].FLOATBUF0\[16\].TE_B
+ VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z sky130_fd_sc_hd__ebufn_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[1\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CLKINV_88 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__inv_1
XFILLER_89_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_57_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_44_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_12_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_60_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CG net13 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[3\] Do0_REG.CLKBUF\[4\] BYTE\[4\].FLOATBUF0\[35\].Z
+ VGND VGND VPWR VPWR Do0[35] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_131_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.DEC0.AND5 SLICE\[3\].RAM8.DEC0.A_buf\[1\] SLICE\[3\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[5\].W.SEL0 sky130_fd_sc_hd__and4b_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_9_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_126_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV_90 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__inv_1
XFILLER_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_67_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_91_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CLKINV_64 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__inv_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_129_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG net117 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CLKINV_173 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__inv_1
XFILLER_10_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_123_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_104_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_106_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_66_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG net73 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_73_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_26_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XEN0BUF.__cell__ EN0 VGND VGND VPWR VPWR DEC0.EN sky130_fd_sc_hd__clkbuf_2
XFILLER_114_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_110_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_63_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG net230 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[7\] Do0_REG.CLKBUF\[0\] BYTE\[0\].FLOATBUF0\[7\].Z
+ VGND VGND VPWR VPWR Do0[7] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_101_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_98_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_74_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_55_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_73_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XDIBUF\[26\].__cell__ Di0[26] VGND VGND VPWR VPWR DIBUF\[26\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG net177 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_123_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_122_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.genblk1.CG net24 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_52_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.genblk1.CLKINV_96 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__inv_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_20_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_109_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[0\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_78_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_65_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_56_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_25_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_24_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_24_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_20_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_79_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV_113 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__inv_1
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG net128 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTIE0\[1\].__cell__ VGND VGND VPWR VPWR TIE0\[1\].__cell__/HI BYTE\[1\].FLOATBUF0\[10\].A
+ sky130_fd_sc_hd__conb_1
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XBYTE\[5\].FLOATBUF0\[44\].__cell__ BYTE\[5\].FLOATBUF0\[40\].A BYTE\[5\].FLOATBUF0\[40\].TE_B
+ VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[0\] Do0_REG.CLKBUF\[1\] BYTE\[1\].FLOATBUF0\[8\].Z
+ VGND VGND VPWR VPWR Do0[8] sky130_fd_sc_hd__dfxtp_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_93_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG net84 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[1\].FLOATBUF0\[12\].__cell__ BYTE\[1\].FLOATBUF0\[10\].A BYTE\[1\].FLOATBUF0\[10\].TE_B
+ VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_61_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_9_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_130_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_97_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_25_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XWEBUF\[6\].__cell__ WE0[6] VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[6\].A sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_121_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_95_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV_145 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__inv_1
XFILLER_31_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[7\] Do0_REG.CLKBUF\[5\] BYTE\[5\].FLOATBUF0\[47\].Z
+ VGND VGND VPWR VPWR Do0[47] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG net197 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_117_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CLKINV_175 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__inv_1
XFILLER_7_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_98_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_93_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_100_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG net188 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.DEC0.AND6 SLICE\[3\].RAM8.DEC0.A_buf\[0\] SLICE\[3\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[6\].W.SEL0 sky130_fd_sc_hd__and4b_2
XFILLER_13_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_8_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_50_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_89_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_66_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDIBUF\[16\].__cell__ Di0[16] VGND VGND VPWR VPWR DIBUF\[16\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_82_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV_211 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__inv_1
XFILLER_5_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_99_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_1_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XDIBUF\[55\].__cell__ Di0[55] VGND VGND VPWR VPWR DIBUF\[55\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_83_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.genblk1.CLKINV_6 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__inv_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_86_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG net95 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_108_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_109_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_2_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XDo0_REG.OUTREG_BYTE\[6\].Do_FF\[0\] Do0_REG.CLKBUF\[6\] BYTE\[6\].FLOATBUF0\[48\].Z
+ VGND VGND VPWR VPWR Do0[48] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_65_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_127_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV_115 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__inv_1
XFILLER_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG net208 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_118_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG net42 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_28_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[32\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_42_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_46_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.Do_CLKBUF\[2\] Do0_REG.CLK_buf VGND VGND VPWR VPWR Do0_REG.CLKBUF\[2\] sky130_fd_sc_hd__clkbuf_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_61_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_68_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG net155 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_84_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_118_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV_147 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__inv_1
XFILLER_106_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[21\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[7\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFBUFENBUF0\[1\].__cell__ EN0 VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[10\].TE_B sky130_fd_sc_hd__clkbuf_2
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_74_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[4\] Do0_REG.CLKBUF\[2\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VGND VGND VPWR VPWR Do0[20] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_90_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_90_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[4\].FLOATBUF0\[36\].__cell__ BYTE\[4\].FLOATBUF0\[32\].A BYTE\[4\].FLOATBUF0\[32\].TE_B
+ VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[36\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_96_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_40_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_109_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_75_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WEBUF\[4\].__cell__ SLICE\[0\].RAM8.WEBUF\[4\].A VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WEBUF\[4\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_98_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_94_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_53_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_61_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_131_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CLKINV_213 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__inv_1
XFILLER_131_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_72_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.DEC0.AND7 SLICE\[3\].RAM8.DEC0.A_buf\[0\] SLICE\[3\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WORD\[7\].W.SEL0 sky130_fd_sc_hd__and4_2
XFILLER_80_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.DEC0.AND0 SLICE\[1\].RAM8.DEC0.A_buf\[0\] SLICE\[1\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[0\].W.SEL0 sky130_fd_sc_hd__nor4b_2
XFILLER_4_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CG net53 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDIBUF\[45\].__cell__ Di0[45] VGND VGND VPWR VPWR DIBUF\[45\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_48_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_129_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WEBUF\[6\].__cell__ SLICE\[0\].RAM8.WEBUF\[6\].A VGND VGND VPWR VPWR
+ SLICE\[2\].RAM8.WEBUF\[6\].X sky130_fd_sc_hd__clkbuf_2
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG net9 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_112_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_1_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG net166 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_73_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.genblk1.CLKINV_117 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__inv_1
XFILLER_41_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_122_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[7\].genblk1.STORAGE DIBUF\[39\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_24_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_117_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV_17 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__inv_1
XFILLER_99_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_113_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_94_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[7\].Do_FF\[4\] Do0_REG.CLKBUF\[7\] BYTE\[7\].FLOATBUF0\[60\].Z
+ VGND VGND VPWR VPWR Do0[60] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG net113 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_10_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_2_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_2_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_127_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CLKINV_149 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_96_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[6\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG net226 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_59_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_86_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_28_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[17\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_11_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_124_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_105_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.DEC0.ABUF\[0\] A0BUF\[0\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.DEC0.A_buf\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.genblk1.CG net64 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_123_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_106_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[6\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG net20 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_90_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_70_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_99_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[7\].genblk1.STORAGE DIBUF\[47\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_97_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].genblk1.STORAGE DIBUF\[59\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CLKINV_215 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__inv_1
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_61_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XBYTE\[3\].FLOATBUF0\[28\].__cell__ BYTE\[3\].FLOATBUF0\[24\].A BYTE\[3\].FLOATBUF0\[24\].TE_B
+ VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z sky130_fd_sc_hd__ebufn_2
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV_242 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_84_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG net133 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_100_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XDIBUF\[35\].__cell__ Di0[35] VGND VGND VPWR VPWR DIBUF\[35\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_75_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_71_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG net124 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_8_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[62\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.genblk1.CLKINV_13 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__inv_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[7\].genblk1.STORAGE DIBUF\[55\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_62_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV_25 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__inv_1
XBYTE\[6\].FLOATBUF0\[51\].__cell__ BYTE\[6\].FLOATBUF0\[48\].A BYTE\[6\].FLOATBUF0\[48\].TE_B
+ VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[51\].Z sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].genblk1.STORAGE DIBUF\[38\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.genblk1.CLKINV_119 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__inv_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[2\].genblk1.STORAGE DIBUF\[50\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[1\].genblk1.STORAGE DIBUF\[33\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_37_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_107_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.DEC0.AND1 SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[0\] SLICE\[1\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[1\].W.SEL0 sky130_fd_sc_hd__and4bb_2
XFILLER_5_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_96_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG net237 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_76_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_117_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[4\].Do_FF\[1\] Do0_REG.CLKBUF\[4\] BYTE\[4\].FLOATBUF0\[33\].Z
+ VGND VGND VPWR VPWR Do0[33] sky130_fd_sc_hd__dfxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG net193 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_39_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_22_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_41_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_103_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_82_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV_178 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[1\].genblk1.STORAGE DIBUF\[41\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_5_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_126_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.genblk1.CG net31 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_76_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[5\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_99_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_117_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_132_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_2_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.genblk1.CG net144 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_60_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.genblk1.CLKINV_8 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__inv_1
XFILLER_9_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].genblk1.STORAGE DIBUF\[63\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[6\].genblk1.STORAGE DIBUF\[46\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_36_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[2\].genblk1.STORAGE DIBUF\[58\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[5\] Do0_REG.CLKBUF\[0\] BYTE\[0\].FLOATBUF0\[5\].Z
+ VGND VGND VPWR VPWR Do0[5] sky130_fd_sc_hd__dfxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_86_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_74_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[2\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[7\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_70_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG net91 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_2_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV_244 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__inv_1
XFILLER_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_46_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_61_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[4\].B.genblk1.CLKINV_21 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__inv_1
XFILLER_127_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_96_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV_33 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__inv_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CG net248 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_110_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_64_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_37_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[50\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[6\].genblk1.STORAGE DIBUF\[54\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_106_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XDIBUF\[25\].__cell__ Di0[25] VGND VGND VPWR VPWR DIBUF\[25\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_133_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[29\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_58_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.BIT\[5\].genblk1.STORAGE DIBUF\[37\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[4\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_74_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].genblk1.STORAGE DIBUF\[49\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG net204 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_16_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[0\].genblk1.STORAGE DIBUF\[32\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_130_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_93_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[58\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_88_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[39\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_37_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_71_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[18\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.BIT\[5\].genblk1.STORAGE DIBUF\[45\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[20\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[0\].genblk1.STORAGE DIBUF\[40\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[7\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[47\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_94_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XDIBUF\[9\].__cell__ Di0[9] VGND VGND VPWR VPWR DIBUF\[9\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_54_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[48\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[38\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[6\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTIE0\[0\].__cell__ VGND VGND VPWR VPWR TIE0\[0\].__cell__/HI BYTE\[0\].FLOATBUF0\[0\].A
+ sky130_fd_sc_hd__conb_1
XFILLER_116_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_130_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV_65 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__inv_1
XBYTE\[5\].FLOATBUF0\[43\].__cell__ BYTE\[5\].FLOATBUF0\[40\].A BYTE\[5\].FLOATBUF0\[40\].TE_B
+ VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[1\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[28\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.genblk1.CLKINV_39 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.DEC0.AND2 SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[1\] SLICE\[1\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[2\].W.SEL0 sky130_fd_sc_hd__and4bb_2
XFILLER_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XBYTE\[1\].FLOATBUF0\[11\].__cell__ BYTE\[1\].FLOATBUF0\[10\].A BYTE\[1\].FLOATBUF0\[10\].TE_B
+ VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_122_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_95_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[7\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_48_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_75_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_44_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[19\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_90_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDo0_REG.OUTREG_BYTE\[5\].Do_FF\[5\] Do0_REG.CLKBUF\[5\] BYTE\[5\].FLOATBUF0\[45\].Z
+ VGND VGND VPWR VPWR Do0[45] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_129_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[4\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ sky130_fd_sc_hd__clkbuf_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.genblk1.CG net102 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[5\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_4_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_112_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.BIT\[6\].genblk1.STORAGE DIBUF\[62\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[7\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_66_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XWEBUF\[5\].__cell__ WE0[5] VGND VGND VPWR VPWR SLICE\[0\].RAM8.WEBUF\[5\].A sky130_fd_sc_hd__clkbuf_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[37\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[9\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[1\].genblk1.STORAGE DIBUF\[57\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_104_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_106_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[5\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[5\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_122_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV_131 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__inv_1
XFILLER_13_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.genblk1.CG net215 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG net49 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[1\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[57\].Z
+ sky130_fd_sc_hd__ebufn_2
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV_41 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__inv_1
XFILLER_8_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_133_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_59_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[7\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[63\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.genblk1.CLKINV_246 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__inv_1
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_23_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[26\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_117_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.BIT\[5\].genblk1.STORAGE DIBUF\[53\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[6\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_133_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[4\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[4\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[4\].genblk1.STORAGE DIBUF\[36\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_26_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[0\].genblk1.STORAGE DIBUF\[48\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_41_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG net162 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_115_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[44\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_5_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[0\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[56\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_83_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[46\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_37_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XDIBUF\[15\].__cell__ Di0[15] VGND VGND VPWR VPWR DIBUF\[15\].X sky130_fd_sc_hd__clkbuf_16
XFILLER_114_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[7\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[25\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[15\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_70_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_109_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDIBUF\[54\].__cell__ Di0[54] VGND VGND VPWR VPWR DIBUF\[54\].X sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_10_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_128_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[27\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_109_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_105_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[6\]
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[54\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[45\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[4\].genblk1.STORAGE DIBUF\[44\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_5_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[0\].genblk1.STORAGE DIBUF\[56\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XFILLER_96_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[8\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV_73 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__inv_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[14\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_102_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[7\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_74_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[6\].B.genblk1.CLKINV_47 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__inv_1
XFILLER_15_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_11_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_7_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV_59 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__inv_1
XFILLER_124_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_93_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CG net69 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_78_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.genblk1.CLKINV_101 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__inv_1
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_1__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[16\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDo0_REG.Do_CLKBUF\[0\] Do0_REG.CLK_buf VGND VGND VPWR VPWR Do0_REG.CLKBUF\[0\] sky130_fd_sc_hd__clkbuf_4
XFILLER_34_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[3\]
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[43\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_30_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XFILLER_128_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[34\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG net60 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_52_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.BIT\[5\].genblk1.STORAGE DIBUF\[61\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[7\].B.Q_WIRE\[5\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_119_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.BIT\[3\].genblk1.STORAGE DIBUF\[35\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[4\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_133_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_102_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[24\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[52\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_16_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[2\] Do0_REG.CLKBUF\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VGND VGND VPWR VPWR Do0[18] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[3\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[3\].W.SEL0 VGND VGND VPWR
+ VPWR SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_109_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[5\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_125_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_1__leaf_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFBUFENBUF0\[0\].__cell__ EN0 VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].TE_B sky130_fd_sc_hd__clkbuf_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[23\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.genblk1.CG net173 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[4\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[4\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[33\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[4\].B.genblk1.CLKINV_133 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__inv_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[4\]
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[60\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.BIT\[2\].genblk1.STORAGE DIBUF\[34\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[4\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[5\].B.genblk1.CLKINV_190 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__inv_1
XFILLER_111_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[11\].Z
+ sky130_fd_sc_hd__ebufn_2
XBYTE\[4\].FLOATBUF0\[35\].__cell__ BYTE\[4\].FLOATBUF0\[32\].A BYTE\[4\].FLOATBUF0\[32\].TE_B
+ VGND VGND VPWR VPWR BYTE\[4\].FLOATBUF0\[35\].Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[13\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.DEC0.AND3 SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[0\] SLICE\[1\].RAM8.DEC0.EN_buf VGND VGND VPWR VPWR
+ SLICE\[1\].RAM8.WORD\[3\].W.SEL0 sky130_fd_sc_hd__and4b_2
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE
+ sky130_fd_sc_hd__and2_1
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG net129 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[53\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X clknet_1_1__leaf_SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XFILLER_91_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV_218 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__inv_1
XFILLER_91_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.genblk1.CLKINV_79 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__inv_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.BIT\[3\].genblk1.STORAGE DIBUF\[43\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[5\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.BIT\[4\].genblk1.STORAGE DIBUF\[52\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X clknet_1_0__leaf_SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[4\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[7\].B.genblk1.CLKINV_248 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__inv_1
XFILLER_31_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\]
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[31\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[4\].B.SEL0_B sky130_fd_sc_hd__inv_1
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[41\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_113_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XFILLER_113_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[2\].FLOATBUF0\[22\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XSLICE\[2\].RAM8.DEC0.ABUF\[1\] A0BUF\[1\].X VGND VGND VPWR VPWR SLICE\[2\].RAM8.DEC0.A_buf\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B sky130_fd_sc_hd__inv_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.Q_WIRE\[3\]
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[59\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[3\].RAM8.WEBUF\[3\].__cell__ SLICE\[0\].RAM8.WEBUF\[3\].A VGND VGND VPWR VPWR
+ SLICE\[3\].RAM8.WEBUF\[3\].X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.Q_WIRE\[5\]
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[7\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[7\].FLOATBUF0\[61\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] sky130_fd_sc_hd__dlxtp_1
XFILLER_58_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X clknet_1_0__leaf_SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] sky130_fd_sc_hd__dlxtp_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\]
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[1\].FLOATBUF0\[12\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[6\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.Q_WIRE\[1\]
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[6\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[6\].FLOATBUF0\[49\].Z
+ sky130_fd_sc_hd__ebufn_2
Xclkbuf_1_0__f_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK clknet_0_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR clknet_1_0__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ sky130_fd_sc_hd__clkbuf_16
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.BIT\[3\].genblk1.STORAGE DIBUF\[51\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[6\].B.Q_WIRE\[3\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.BIT\[2\].genblk1.STORAGE DIBUF\[42\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[5\].B.Q_WIRE\[2\] sky130_fd_sc_hd__dlxtp_1
XFILLER_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[0\].FLOATBUF0\[0\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X clknet_1_0__leaf_SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] sky130_fd_sc_hd__dlxtp_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\]
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[3\].FLOATBUF0\[30\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_91_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.Q_WIRE\[0\]
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[40\].Z
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.Q_WIRE\[2\]
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[5\].B.SEL0_B VGND VGND VPWR VPWR BYTE\[5\].FLOATBUF0\[42\].Z
+ sky130_fd_sc_hd__ebufn_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG net233 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE
+ VGND VGND VPWR VPWR SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK sky130_fd_sc_hd__dlclkp_1
XFILLER_118_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.BIT\[4\].genblk1.STORAGE DIBUF\[60\].X clknet_1_1__leaf_SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.GCLK
+ VGND VGND VPWR VPWR SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[7\].B.Q_WIRE\[4\] sky130_fd_sc_hd__dlxtp_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ VGND VGND VPWR VPWR clknet_0_SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

