module logo();
endmodule
