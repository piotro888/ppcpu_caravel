magic
tech sky130B
magscale 1 2
timestamp 1662672544
<< obsli1 >>
rect 1104 2159 170752 171377
<< obsm1 >>
rect 14 1708 171382 171408
<< metal2 >>
rect 1950 173277 2006 174077
rect 6458 173277 6514 174077
rect 10322 173277 10378 174077
rect 14186 173277 14242 174077
rect 18050 173277 18106 174077
rect 21914 173277 21970 174077
rect 25778 173277 25834 174077
rect 29642 173277 29698 174077
rect 33506 173277 33562 174077
rect 37370 173277 37426 174077
rect 41234 173277 41290 174077
rect 45098 173277 45154 174077
rect 48962 173277 49018 174077
rect 52826 173277 52882 174077
rect 56690 173277 56746 174077
rect 60554 173277 60610 174077
rect 64418 173277 64474 174077
rect 68282 173277 68338 174077
rect 72146 173277 72202 174077
rect 76010 173277 76066 174077
rect 79874 173277 79930 174077
rect 83738 173277 83794 174077
rect 88246 173277 88302 174077
rect 92110 173277 92166 174077
rect 95974 173277 96030 174077
rect 99838 173277 99894 174077
rect 103702 173277 103758 174077
rect 107566 173277 107622 174077
rect 111430 173277 111486 174077
rect 115294 173277 115350 174077
rect 119158 173277 119214 174077
rect 123022 173277 123078 174077
rect 126886 173277 126942 174077
rect 130750 173277 130806 174077
rect 134614 173277 134670 174077
rect 138478 173277 138534 174077
rect 142342 173277 142398 174077
rect 146206 173277 146262 174077
rect 150070 173277 150126 174077
rect 153934 173277 153990 174077
rect 157798 173277 157854 174077
rect 161662 173277 161718 174077
rect 165526 173277 165582 174077
rect 169390 173277 169446 174077
rect 18 0 74 800
rect 3882 0 3938 800
rect 7746 0 7802 800
rect 11610 0 11666 800
rect 15474 0 15530 800
rect 19338 0 19394 800
rect 23202 0 23258 800
rect 27066 0 27122 800
rect 30930 0 30986 800
rect 34794 0 34850 800
rect 38658 0 38714 800
rect 42522 0 42578 800
rect 46386 0 46442 800
rect 50250 0 50306 800
rect 54114 0 54170 800
rect 57978 0 58034 800
rect 61842 0 61898 800
rect 65706 0 65762 800
rect 69570 0 69626 800
rect 73434 0 73490 800
rect 77298 0 77354 800
rect 81162 0 81218 800
rect 85670 0 85726 800
rect 89534 0 89590 800
rect 93398 0 93454 800
rect 97262 0 97318 800
rect 101126 0 101182 800
rect 104990 0 105046 800
rect 108854 0 108910 800
rect 112718 0 112774 800
rect 116582 0 116638 800
rect 120446 0 120502 800
rect 124310 0 124366 800
rect 128174 0 128230 800
rect 132038 0 132094 800
rect 135902 0 135958 800
rect 139766 0 139822 800
rect 143630 0 143686 800
rect 147494 0 147550 800
rect 151358 0 151414 800
rect 155222 0 155278 800
rect 159086 0 159142 800
rect 162950 0 163006 800
rect 166814 0 166870 800
rect 171322 0 171378 800
<< obsm2 >>
rect 20 173221 1894 173277
rect 2062 173221 6402 173277
rect 6570 173221 10266 173277
rect 10434 173221 14130 173277
rect 14298 173221 17994 173277
rect 18162 173221 21858 173277
rect 22026 173221 25722 173277
rect 25890 173221 29586 173277
rect 29754 173221 33450 173277
rect 33618 173221 37314 173277
rect 37482 173221 41178 173277
rect 41346 173221 45042 173277
rect 45210 173221 48906 173277
rect 49074 173221 52770 173277
rect 52938 173221 56634 173277
rect 56802 173221 60498 173277
rect 60666 173221 64362 173277
rect 64530 173221 68226 173277
rect 68394 173221 72090 173277
rect 72258 173221 75954 173277
rect 76122 173221 79818 173277
rect 79986 173221 83682 173277
rect 83850 173221 88190 173277
rect 88358 173221 92054 173277
rect 92222 173221 95918 173277
rect 96086 173221 99782 173277
rect 99950 173221 103646 173277
rect 103814 173221 107510 173277
rect 107678 173221 111374 173277
rect 111542 173221 115238 173277
rect 115406 173221 119102 173277
rect 119270 173221 122966 173277
rect 123134 173221 126830 173277
rect 126998 173221 130694 173277
rect 130862 173221 134558 173277
rect 134726 173221 138422 173277
rect 138590 173221 142286 173277
rect 142454 173221 146150 173277
rect 146318 173221 150014 173277
rect 150182 173221 153878 173277
rect 154046 173221 157742 173277
rect 157910 173221 161606 173277
rect 161774 173221 165470 173277
rect 165638 173221 169334 173277
rect 169502 173221 171376 173277
rect 20 856 171376 173221
rect 130 800 3826 856
rect 3994 800 7690 856
rect 7858 800 11554 856
rect 11722 800 15418 856
rect 15586 800 19282 856
rect 19450 800 23146 856
rect 23314 800 27010 856
rect 27178 800 30874 856
rect 31042 800 34738 856
rect 34906 800 38602 856
rect 38770 800 42466 856
rect 42634 800 46330 856
rect 46498 800 50194 856
rect 50362 800 54058 856
rect 54226 800 57922 856
rect 58090 800 61786 856
rect 61954 800 65650 856
rect 65818 800 69514 856
rect 69682 800 73378 856
rect 73546 800 77242 856
rect 77410 800 81106 856
rect 81274 800 85614 856
rect 85782 800 89478 856
rect 89646 800 93342 856
rect 93510 800 97206 856
rect 97374 800 101070 856
rect 101238 800 104934 856
rect 105102 800 108798 856
rect 108966 800 112662 856
rect 112830 800 116526 856
rect 116694 800 120390 856
rect 120558 800 124254 856
rect 124422 800 128118 856
rect 128286 800 131982 856
rect 132150 800 135846 856
rect 136014 800 139710 856
rect 139878 800 143574 856
rect 143742 800 147438 856
rect 147606 800 151302 856
rect 151470 800 155166 856
rect 155334 800 159030 856
rect 159198 800 162894 856
rect 163062 800 166758 856
rect 166926 800 171266 856
<< metal3 >>
rect 0 172048 800 172168
rect 171133 171368 171933 171488
rect 0 167968 800 168088
rect 171133 167288 171933 167408
rect 0 163888 800 164008
rect 171133 163208 171933 163328
rect 0 159808 800 159928
rect 171133 159128 171933 159248
rect 0 155728 800 155848
rect 171133 155048 171933 155168
rect 0 151648 800 151768
rect 171133 150968 171933 151088
rect 0 147568 800 147688
rect 171133 146888 171933 147008
rect 0 143488 800 143608
rect 171133 142808 171933 142928
rect 0 139408 800 139528
rect 171133 138728 171933 138848
rect 0 135328 800 135448
rect 171133 134648 171933 134768
rect 0 131248 800 131368
rect 171133 130568 171933 130688
rect 0 127168 800 127288
rect 171133 126488 171933 126608
rect 0 123088 800 123208
rect 171133 122408 171933 122528
rect 0 119008 800 119128
rect 171133 118328 171933 118448
rect 0 114928 800 115048
rect 171133 114248 171933 114368
rect 0 110848 800 110968
rect 171133 110168 171933 110288
rect 0 106768 800 106888
rect 171133 106088 171933 106208
rect 0 102688 800 102808
rect 171133 102008 171933 102128
rect 0 98608 800 98728
rect 171133 97928 171933 98048
rect 0 94528 800 94648
rect 171133 93848 171933 93968
rect 0 90448 800 90568
rect 171133 89768 171933 89888
rect 0 85688 800 85808
rect 171133 85688 171933 85808
rect 0 81608 800 81728
rect 171133 80928 171933 81048
rect 0 77528 800 77648
rect 171133 76848 171933 76968
rect 0 73448 800 73568
rect 171133 72768 171933 72888
rect 0 69368 800 69488
rect 171133 68688 171933 68808
rect 0 65288 800 65408
rect 171133 64608 171933 64728
rect 0 61208 800 61328
rect 171133 60528 171933 60648
rect 0 57128 800 57248
rect 171133 56448 171933 56568
rect 0 53048 800 53168
rect 171133 52368 171933 52488
rect 0 48968 800 49088
rect 171133 48288 171933 48408
rect 0 44888 800 45008
rect 171133 44208 171933 44328
rect 0 40808 800 40928
rect 171133 40128 171933 40248
rect 0 36728 800 36848
rect 171133 36048 171933 36168
rect 0 32648 800 32768
rect 171133 31968 171933 32088
rect 0 28568 800 28688
rect 171133 27888 171933 28008
rect 0 24488 800 24608
rect 171133 23808 171933 23928
rect 0 20408 800 20528
rect 171133 19728 171933 19848
rect 0 16328 800 16448
rect 171133 15648 171933 15768
rect 0 12248 800 12368
rect 171133 11568 171933 11688
rect 0 8168 800 8288
rect 171133 7488 171933 7608
rect 0 4088 800 4208
rect 171133 3408 171933 3528
<< obsm3 >>
rect 880 171968 171133 172141
rect 800 171568 171133 171968
rect 800 171288 171053 171568
rect 800 168168 171133 171288
rect 880 167888 171133 168168
rect 800 167488 171133 167888
rect 800 167208 171053 167488
rect 800 164088 171133 167208
rect 880 163808 171133 164088
rect 800 163408 171133 163808
rect 800 163128 171053 163408
rect 800 160008 171133 163128
rect 880 159728 171133 160008
rect 800 159328 171133 159728
rect 800 159048 171053 159328
rect 800 155928 171133 159048
rect 880 155648 171133 155928
rect 800 155248 171133 155648
rect 800 154968 171053 155248
rect 800 151848 171133 154968
rect 880 151568 171133 151848
rect 800 151168 171133 151568
rect 800 150888 171053 151168
rect 800 147768 171133 150888
rect 880 147488 171133 147768
rect 800 147088 171133 147488
rect 800 146808 171053 147088
rect 800 143688 171133 146808
rect 880 143408 171133 143688
rect 800 143008 171133 143408
rect 800 142728 171053 143008
rect 800 139608 171133 142728
rect 880 139328 171133 139608
rect 800 138928 171133 139328
rect 800 138648 171053 138928
rect 800 135528 171133 138648
rect 880 135248 171133 135528
rect 800 134848 171133 135248
rect 800 134568 171053 134848
rect 800 131448 171133 134568
rect 880 131168 171133 131448
rect 800 130768 171133 131168
rect 800 130488 171053 130768
rect 800 127368 171133 130488
rect 880 127088 171133 127368
rect 800 126688 171133 127088
rect 800 126408 171053 126688
rect 800 123288 171133 126408
rect 880 123008 171133 123288
rect 800 122608 171133 123008
rect 800 122328 171053 122608
rect 800 119208 171133 122328
rect 880 118928 171133 119208
rect 800 118528 171133 118928
rect 800 118248 171053 118528
rect 800 115128 171133 118248
rect 880 114848 171133 115128
rect 800 114448 171133 114848
rect 800 114168 171053 114448
rect 800 111048 171133 114168
rect 880 110768 171133 111048
rect 800 110368 171133 110768
rect 800 110088 171053 110368
rect 800 106968 171133 110088
rect 880 106688 171133 106968
rect 800 106288 171133 106688
rect 800 106008 171053 106288
rect 800 102888 171133 106008
rect 880 102608 171133 102888
rect 800 102208 171133 102608
rect 800 101928 171053 102208
rect 800 98808 171133 101928
rect 880 98528 171133 98808
rect 800 98128 171133 98528
rect 800 97848 171053 98128
rect 800 94728 171133 97848
rect 880 94448 171133 94728
rect 800 94048 171133 94448
rect 800 93768 171053 94048
rect 800 90648 171133 93768
rect 880 90368 171133 90648
rect 800 89968 171133 90368
rect 800 89688 171053 89968
rect 800 85888 171133 89688
rect 880 85608 171053 85888
rect 800 81808 171133 85608
rect 880 81528 171133 81808
rect 800 81128 171133 81528
rect 800 80848 171053 81128
rect 800 77728 171133 80848
rect 880 77448 171133 77728
rect 800 77048 171133 77448
rect 800 76768 171053 77048
rect 800 73648 171133 76768
rect 880 73368 171133 73648
rect 800 72968 171133 73368
rect 800 72688 171053 72968
rect 800 69568 171133 72688
rect 880 69288 171133 69568
rect 800 68888 171133 69288
rect 800 68608 171053 68888
rect 800 65488 171133 68608
rect 880 65208 171133 65488
rect 800 64808 171133 65208
rect 800 64528 171053 64808
rect 800 61408 171133 64528
rect 880 61128 171133 61408
rect 800 60728 171133 61128
rect 800 60448 171053 60728
rect 800 57328 171133 60448
rect 880 57048 171133 57328
rect 800 56648 171133 57048
rect 800 56368 171053 56648
rect 800 53248 171133 56368
rect 880 52968 171133 53248
rect 800 52568 171133 52968
rect 800 52288 171053 52568
rect 800 49168 171133 52288
rect 880 48888 171133 49168
rect 800 48488 171133 48888
rect 800 48208 171053 48488
rect 800 45088 171133 48208
rect 880 44808 171133 45088
rect 800 44408 171133 44808
rect 800 44128 171053 44408
rect 800 41008 171133 44128
rect 880 40728 171133 41008
rect 800 40328 171133 40728
rect 800 40048 171053 40328
rect 800 36928 171133 40048
rect 880 36648 171133 36928
rect 800 36248 171133 36648
rect 800 35968 171053 36248
rect 800 32848 171133 35968
rect 880 32568 171133 32848
rect 800 32168 171133 32568
rect 800 31888 171053 32168
rect 800 28768 171133 31888
rect 880 28488 171133 28768
rect 800 28088 171133 28488
rect 800 27808 171053 28088
rect 800 24688 171133 27808
rect 880 24408 171133 24688
rect 800 24008 171133 24408
rect 800 23728 171053 24008
rect 800 20608 171133 23728
rect 880 20328 171133 20608
rect 800 19928 171133 20328
rect 800 19648 171053 19928
rect 800 16528 171133 19648
rect 880 16248 171133 16528
rect 800 15848 171133 16248
rect 800 15568 171053 15848
rect 800 12448 171133 15568
rect 880 12168 171133 12448
rect 800 11768 171133 12168
rect 800 11488 171053 11768
rect 800 8368 171133 11488
rect 880 8088 171133 8368
rect 800 7688 171133 8088
rect 800 7408 171053 7688
rect 800 4288 171133 7408
rect 880 4008 171133 4288
rect 800 3608 171133 4008
rect 800 3328 171053 3608
rect 800 2143 171133 3328
<< metal4 >>
rect 4208 2128 4528 171408
rect 19568 2128 19888 171408
rect 34928 2128 35248 171408
rect 50288 2128 50608 171408
rect 65648 2128 65968 171408
rect 81008 2128 81328 171408
rect 96368 2128 96688 171408
rect 111728 2128 112048 171408
rect 127088 2128 127408 171408
rect 142448 2128 142768 171408
rect 157808 2128 158128 171408
<< obsm4 >>
rect 2267 171488 169405 171733
rect 2267 2347 4128 171488
rect 4608 2347 19488 171488
rect 19968 2347 34848 171488
rect 35328 2347 50208 171488
rect 50688 2347 65568 171488
rect 66048 2347 80928 171488
rect 81408 2347 96288 171488
rect 96768 2347 111648 171488
rect 112128 2347 127008 171488
rect 127488 2347 142368 171488
rect 142848 2347 157728 171488
rect 158208 2347 169405 171488
<< metal5 >>
rect 1056 158526 170800 158846
rect 1056 143208 170800 143528
rect 1056 127890 170800 128210
rect 1056 112572 170800 112892
rect 1056 97254 170800 97574
rect 1056 81936 170800 82256
rect 1056 66618 170800 66938
rect 1056 51300 170800 51620
rect 1056 35982 170800 36302
rect 1056 20664 170800 20984
rect 1056 5346 170800 5666
<< labels >>
rlabel metal4 s 19568 2128 19888 171408 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 171408 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 171408 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 171408 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 171408 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 20664 170800 20984 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 51300 170800 51620 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 81936 170800 82256 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 112572 170800 112892 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 143208 170800 143528 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 171408 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 171408 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 171408 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 171408 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 171408 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 171408 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 170800 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 170800 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66618 170800 66938 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 97254 170800 97574 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 127890 170800 128210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 158526 170800 158846 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 165526 173277 165582 174077 6 i_addr[0]
port 3 nsew signal input
rlabel metal2 s 68282 173277 68338 174077 6 i_addr[1]
port 4 nsew signal input
rlabel metal3 s 171133 23808 171933 23928 6 i_addr[2]
port 5 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 i_addr[3]
port 6 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 i_addr[4]
port 7 nsew signal input
rlabel metal2 s 21914 173277 21970 174077 6 i_addr[5]
port 8 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 i_clk
port 9 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 i_data[0]
port 10 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 i_data[10]
port 11 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 i_data[11]
port 12 nsew signal input
rlabel metal3 s 171133 163208 171933 163328 6 i_data[12]
port 13 nsew signal input
rlabel metal2 s 111430 173277 111486 174077 6 i_data[13]
port 14 nsew signal input
rlabel metal2 s 103702 173277 103758 174077 6 i_data[14]
port 15 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 i_data[15]
port 16 nsew signal input
rlabel metal2 s 79874 173277 79930 174077 6 i_data[16]
port 17 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 i_data[17]
port 18 nsew signal input
rlabel metal2 s 14186 173277 14242 174077 6 i_data[18]
port 19 nsew signal input
rlabel metal3 s 0 172048 800 172168 6 i_data[19]
port 20 nsew signal input
rlabel metal2 s 99838 173277 99894 174077 6 i_data[1]
port 21 nsew signal input
rlabel metal3 s 171133 27888 171933 28008 6 i_data[20]
port 22 nsew signal input
rlabel metal2 s 37370 173277 37426 174077 6 i_data[21]
port 23 nsew signal input
rlabel metal2 s 76010 173277 76066 174077 6 i_data[22]
port 24 nsew signal input
rlabel metal3 s 171133 76848 171933 76968 6 i_data[23]
port 25 nsew signal input
rlabel metal2 s 41234 173277 41290 174077 6 i_data[24]
port 26 nsew signal input
rlabel metal3 s 171133 155048 171933 155168 6 i_data[25]
port 27 nsew signal input
rlabel metal3 s 171133 15648 171933 15768 6 i_data[26]
port 28 nsew signal input
rlabel metal2 s 130750 173277 130806 174077 6 i_data[27]
port 29 nsew signal input
rlabel metal3 s 171133 11568 171933 11688 6 i_data[28]
port 30 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 i_data[29]
port 31 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 i_data[2]
port 32 nsew signal input
rlabel metal2 s 10322 173277 10378 174077 6 i_data[30]
port 33 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 i_data[31]
port 34 nsew signal input
rlabel metal3 s 171133 146888 171933 147008 6 i_data[32]
port 35 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 i_data[33]
port 36 nsew signal input
rlabel metal2 s 33506 173277 33562 174077 6 i_data[34]
port 37 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 i_data[35]
port 38 nsew signal input
rlabel metal2 s 153934 173277 153990 174077 6 i_data[36]
port 39 nsew signal input
rlabel metal2 s 6458 173277 6514 174077 6 i_data[37]
port 40 nsew signal input
rlabel metal2 s 52826 173277 52882 174077 6 i_data[38]
port 41 nsew signal input
rlabel metal3 s 171133 138728 171933 138848 6 i_data[39]
port 42 nsew signal input
rlabel metal3 s 171133 110168 171933 110288 6 i_data[3]
port 43 nsew signal input
rlabel metal3 s 171133 72768 171933 72888 6 i_data[40]
port 44 nsew signal input
rlabel metal2 s 138478 173277 138534 174077 6 i_data[41]
port 45 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 i_data[42]
port 46 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 i_data[43]
port 47 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 i_data[44]
port 48 nsew signal input
rlabel metal3 s 171133 134648 171933 134768 6 i_data[45]
port 49 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 i_data[46]
port 50 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 i_data[47]
port 51 nsew signal input
rlabel metal3 s 171133 93848 171933 93968 6 i_data[48]
port 52 nsew signal input
rlabel metal2 s 161662 173277 161718 174077 6 i_data[49]
port 53 nsew signal input
rlabel metal2 s 72146 173277 72202 174077 6 i_data[4]
port 54 nsew signal input
rlabel metal3 s 171133 85688 171933 85808 6 i_data[50]
port 55 nsew signal input
rlabel metal2 s 157798 173277 157854 174077 6 i_data[51]
port 56 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 i_data[52]
port 57 nsew signal input
rlabel metal3 s 171133 36048 171933 36168 6 i_data[53]
port 58 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 i_data[54]
port 59 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 i_data[55]
port 60 nsew signal input
rlabel metal2 s 150070 173277 150126 174077 6 i_data[56]
port 61 nsew signal input
rlabel metal3 s 171133 171368 171933 171488 6 i_data[57]
port 62 nsew signal input
rlabel metal2 s 64418 173277 64474 174077 6 i_data[58]
port 63 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 i_data[59]
port 64 nsew signal input
rlabel metal2 s 107566 173277 107622 174077 6 i_data[5]
port 65 nsew signal input
rlabel metal2 s 18050 173277 18106 174077 6 i_data[60]
port 66 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 i_data[61]
port 67 nsew signal input
rlabel metal3 s 0 167968 800 168088 6 i_data[62]
port 68 nsew signal input
rlabel metal3 s 0 151648 800 151768 6 i_data[63]
port 69 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 i_data[64]
port 70 nsew signal input
rlabel metal2 s 146206 173277 146262 174077 6 i_data[65]
port 71 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 i_data[66]
port 72 nsew signal input
rlabel metal3 s 171133 44208 171933 44328 6 i_data[67]
port 73 nsew signal input
rlabel metal3 s 171133 64608 171933 64728 6 i_data[68]
port 74 nsew signal input
rlabel metal3 s 0 163888 800 164008 6 i_data[69]
port 75 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 i_data[6]
port 76 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 i_data[70]
port 77 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 i_data[71]
port 78 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 i_data[72]
port 79 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 i_data[73]
port 80 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 i_data[74]
port 81 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 i_data[75]
port 82 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 i_data[76]
port 83 nsew signal input
rlabel metal2 s 48962 173277 49018 174077 6 i_data[77]
port 84 nsew signal input
rlabel metal2 s 60554 173277 60610 174077 6 i_data[78]
port 85 nsew signal input
rlabel metal3 s 0 131248 800 131368 6 i_data[79]
port 86 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 i_data[7]
port 87 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 i_data[80]
port 88 nsew signal input
rlabel metal3 s 171133 142808 171933 142928 6 i_data[81]
port 89 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 i_data[8]
port 90 nsew signal input
rlabel metal3 s 0 155728 800 155848 6 i_data[9]
port 91 nsew signal input
rlabel metal3 s 171133 122408 171933 122528 6 i_rst
port 92 nsew signal input
rlabel metal2 s 45098 173277 45154 174077 6 i_we
port 93 nsew signal input
rlabel metal3 s 171133 48288 171933 48408 6 o_data[0]
port 94 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 o_data[10]
port 95 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 o_data[11]
port 96 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 o_data[12]
port 97 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 o_data[13]
port 98 nsew signal output
rlabel metal3 s 171133 89768 171933 89888 6 o_data[14]
port 99 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 o_data[15]
port 100 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 o_data[16]
port 101 nsew signal output
rlabel metal2 s 92110 173277 92166 174077 6 o_data[17]
port 102 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 o_data[18]
port 103 nsew signal output
rlabel metal3 s 0 159808 800 159928 6 o_data[19]
port 104 nsew signal output
rlabel metal3 s 171133 159128 171933 159248 6 o_data[1]
port 105 nsew signal output
rlabel metal3 s 171133 56448 171933 56568 6 o_data[20]
port 106 nsew signal output
rlabel metal2 s 95974 173277 96030 174077 6 o_data[21]
port 107 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 o_data[22]
port 108 nsew signal output
rlabel metal2 s 115294 173277 115350 174077 6 o_data[23]
port 109 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 o_data[24]
port 110 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 o_data[25]
port 111 nsew signal output
rlabel metal3 s 171133 19728 171933 19848 6 o_data[26]
port 112 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 o_data[27]
port 113 nsew signal output
rlabel metal3 s 171133 130568 171933 130688 6 o_data[28]
port 114 nsew signal output
rlabel metal3 s 171133 97928 171933 98048 6 o_data[29]
port 115 nsew signal output
rlabel metal2 s 126886 173277 126942 174077 6 o_data[2]
port 116 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 o_data[30]
port 117 nsew signal output
rlabel metal3 s 171133 40128 171933 40248 6 o_data[31]
port 118 nsew signal output
rlabel metal3 s 171133 102008 171933 102128 6 o_data[32]
port 119 nsew signal output
rlabel metal2 s 56690 173277 56746 174077 6 o_data[33]
port 120 nsew signal output
rlabel metal3 s 171133 68688 171933 68808 6 o_data[34]
port 121 nsew signal output
rlabel metal3 s 171133 3408 171933 3528 6 o_data[35]
port 122 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 o_data[36]
port 123 nsew signal output
rlabel metal3 s 171133 126488 171933 126608 6 o_data[37]
port 124 nsew signal output
rlabel metal2 s 134614 173277 134670 174077 6 o_data[38]
port 125 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 o_data[39]
port 126 nsew signal output
rlabel metal3 s 171133 52368 171933 52488 6 o_data[3]
port 127 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 o_data[40]
port 128 nsew signal output
rlabel metal3 s 171133 7488 171933 7608 6 o_data[41]
port 129 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 o_data[42]
port 130 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 o_data[43]
port 131 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 o_data[44]
port 132 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 o_data[45]
port 133 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 o_data[46]
port 134 nsew signal output
rlabel metal3 s 171133 150968 171933 151088 6 o_data[47]
port 135 nsew signal output
rlabel metal3 s 171133 106088 171933 106208 6 o_data[48]
port 136 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 o_data[49]
port 137 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 o_data[4]
port 138 nsew signal output
rlabel metal3 s 171133 60528 171933 60648 6 o_data[50]
port 139 nsew signal output
rlabel metal3 s 0 114928 800 115048 6 o_data[51]
port 140 nsew signal output
rlabel metal3 s 171133 114248 171933 114368 6 o_data[52]
port 141 nsew signal output
rlabel metal3 s 171133 167288 171933 167408 6 o_data[53]
port 142 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 o_data[54]
port 143 nsew signal output
rlabel metal2 s 169390 173277 169446 174077 6 o_data[55]
port 144 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 o_data[56]
port 145 nsew signal output
rlabel metal3 s 0 127168 800 127288 6 o_data[57]
port 146 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 o_data[58]
port 147 nsew signal output
rlabel metal2 s 18 0 74 800 6 o_data[59]
port 148 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 o_data[5]
port 149 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 o_data[60]
port 150 nsew signal output
rlabel metal2 s 25778 173277 25834 174077 6 o_data[61]
port 151 nsew signal output
rlabel metal2 s 88246 173277 88302 174077 6 o_data[62]
port 152 nsew signal output
rlabel metal3 s 0 110848 800 110968 6 o_data[63]
port 153 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 o_data[64]
port 154 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 o_data[65]
port 155 nsew signal output
rlabel metal2 s 119158 173277 119214 174077 6 o_data[66]
port 156 nsew signal output
rlabel metal2 s 83738 173277 83794 174077 6 o_data[67]
port 157 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 o_data[68]
port 158 nsew signal output
rlabel metal2 s 142342 173277 142398 174077 6 o_data[69]
port 159 nsew signal output
rlabel metal3 s 171133 31968 171933 32088 6 o_data[6]
port 160 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 o_data[70]
port 161 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 o_data[71]
port 162 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 o_data[72]
port 163 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 o_data[73]
port 164 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 o_data[74]
port 165 nsew signal output
rlabel metal3 s 171133 118328 171933 118448 6 o_data[75]
port 166 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 o_data[76]
port 167 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 o_data[77]
port 168 nsew signal output
rlabel metal2 s 123022 173277 123078 174077 6 o_data[78]
port 169 nsew signal output
rlabel metal2 s 1950 173277 2006 174077 6 o_data[79]
port 170 nsew signal output
rlabel metal2 s 29642 173277 29698 174077 6 o_data[7]
port 171 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 o_data[80]
port 172 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 o_data[81]
port 173 nsew signal output
rlabel metal3 s 0 147568 800 147688 6 o_data[8]
port 174 nsew signal output
rlabel metal3 s 171133 80928 171933 81048 6 o_data[9]
port 175 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 171933 174077
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 74645108
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/dffram/runs/22_09_08_23_15/results/signoff/d_dffram.magic.gds
string GDS_START 433096
<< end >>

